VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
	DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

USEMINSPACING OBS ON ;


PROPERTYDEFINITIONS 
END PROPERTYDEFINITIONS
LAYER diff

	TYPE MASTERSLICE ;
END diff

LAYER poly

	TYPE MASTERSLICE ;
END poly

LAYER mcon

	TYPE CUT ;
END mcon

LAYER met1

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.46 ;
	WIDTH 0.14 ;
	OFFSET 0.0 ;
	AREA 0.083 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.14 
		WIDTH 3.0	           		  0.28 ;

	WIREEXTENSION 0.07 ;
	MINWIDTH 0.14 ;
	MINENCLOSEDAREA 0.14 ;
	
	RESISTANCE RPERSQ 0.125 ;
	CAPACITANCE CPERSQDIST 2.57784e-05 ;
	THICKNESS 0.35 ;
	EDGECAPACITANCE 4.0567e-05 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 )  ( 0.0125 400.0 )  ( 0.0225 2609.0 )  ( 22.5 11600.0 ) ) ;
	ACCURRENTDENSITY RMS 6.1 ;
	DCCURRENTDENSITY AVERAGE 2.8 ;
END met1

LAYER via

	TYPE CUT ;
	SPACING 0.17  ;
	
	WIDTH 0.15 ;
	ENCLOSURE  ABOVE  0.055 0.085  ;
	ENCLOSURE  BELOW  0.055 0.085  ;
	
	RESISTANCE 4.5 ;
	DCCURRENTDENSITY AVERAGE 0.29 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 )  ( 0.0125 6.0 )  ( 0.0225 6.81 )  ( 22.5 816.0 ) ) ;
END via

LAYER met2

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.46 ;
	WIDTH 0.14 ;
	OFFSET 0.0 ;
	AREA 0.0676 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.14 
		WIDTH 3.0	           		  0.28 ;

	WIREEXTENSION 0.07 ;
	MINWIDTH 0.14 ;
	MINENCLOSEDAREA 0.14 ;
	
	RESISTANCE RPERSQ 0.125 ;
	CAPACITANCE CPERSQDIST 1.69423e-05 ;
	THICKNESS 0.35 ;
	EDGECAPACITANCE 3.7759e-05 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 )  ( 0.0125 400.0 )  ( 0.0225 2609.0 )  ( 22.5 11600.0 ) ) ;
	ACCURRENTDENSITY RMS 6.1 ;
	DCCURRENTDENSITY AVERAGE 2.8 ;
END met2

LAYER via2

	TYPE CUT ;
	SPACING 0.2  ;
	
	WIDTH 0.2 ;
	ENCLOSURE  ABOVE  0.065 0.065  ;
	ENCLOSURE  BELOW  0.04 0.085  ;
	
	RESISTANCE 3.41 ;
	DCCURRENTDENSITY AVERAGE 0.48 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 )  ( 0.0125 6.0 )  ( 0.0225 6.81 )  ( 22.5 816.0 ) ) ;
END via2

LAYER met3

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 0.69 ;
	WIDTH 0.3 ;
	OFFSET 0.0 ;
	AREA 0.24 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.3 
		WIDTH 3.0	           		  0.4 ;

	WIREEXTENSION 0.15 ;
	MINWIDTH 0.3 ;
	RESISTANCE RPERSQ 0.047 ;
	CAPACITANCE CPERSQDIST 1.23729e-05 ;
	THICKNESS 0.8 ;
	EDGECAPACITANCE 4.0989e-05 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 )  ( 0.0125 400.0 )  ( 0.0225 2609.0 )  ( 22.5 11600.0 ) ) ;
	ACCURRENTDENSITY RMS 14.9 ;
	DCCURRENTDENSITY AVERAGE 6.8 ;
END met3

LAYER via3

	TYPE CUT ;
	SPACING 0.2  ;
	
	WIDTH 0.2 ;
	ENCLOSURE  ABOVE  0.065 0.065  ;
	ENCLOSURE  BELOW  0.06 0.09  ;
	
	RESISTANCE 3.41 ;
	DCCURRENTDENSITY AVERAGE 0.48 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 )  ( 0.0125 6.0 )  ( 0.0225 6.81 )  ( 22.5 816.0 ) ) ;
END via3

LAYER met4

	TYPE ROUTING ;
	DIRECTION VERTICAL ;
	PITCH 0.69 ;
	WIDTH 0.3 ;
	OFFSET 0.0 ;
	AREA 0.24 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  0.3 
		WIDTH 3.0	           		  0.4 ;

	WIREEXTENSION 0.15 ;
	MINWIDTH 0.3 ;
	RESISTANCE RPERSQ 0.047 ;
	CAPACITANCE CPERSQDIST 8.41537e-06 ;
	THICKNESS 0.8 ;
	EDGECAPACITANCE 3.6676e-05 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 )  ( 0.0125 400.0 )  ( 0.0225 2609.0 )  ( 22.5 11600.0 ) ) ;
	ACCURRENTDENSITY RMS 14.9 ;
	DCCURRENTDENSITY AVERAGE 6.8 ;
END met4

LAYER via4

	TYPE CUT ;
	SPACING 0.8  ;
	
	WIDTH 0.8 ;
	ENCLOSURE  ABOVE  0.31 0.31  ;
	ENCLOSURE  BELOW  0.19 0.19  ;
	
	RESISTANCE 0.38 ;
	DCCURRENTDENSITY AVERAGE 2.49 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFAREARATIO PWL ( ( 0.0 6.0 )  ( 0.0125 6.0 )  ( 0.0225 6.81 )  ( 22.5 816.0 ) ) ;
END via4

LAYER met5

	TYPE ROUTING ;
	DIRECTION HORIZONTAL ;
	PITCH 3.22 ;
	WIDTH 1.6 ;
	OFFSET 0.0 ;
	AREA 4.0 ;
	
	SPACINGTABLE  PARALLELRUNLENGTH
		     		 0.0 
		WIDTH 0.0	           		  1.6 ;

	WIREEXTENSION 0.8 ;
	MINWIDTH 1.6 ;
	RESISTANCE RPERSQ 0.029 ;
	CAPACITANCE CPERSQDIST 6.32063e-06 ;
	THICKNESS 1.2 ;
	EDGECAPACITANCE 3.8851e-05 ;
	ANTENNAMODEL OXIDE1 ;
	ANTENNADIFFSIDEAREARATIO PWL ( ( 0.0 400.0 )  ( 0.0125 400.0 )  ( 0.0225 2609.0 )  ( 22.5 11600.0 ) ) ;
	ACCURRENTDENSITY RMS 22.34 ;
	DCCURRENTDENSITY AVERAGE 10.17 ;
END met5

VIARULE M1M2_PR GENERATE 
	LAYER met1 ;
		ENCLOSURE 0.085 0.055 ;
		WIDTH 0 TO 1000 ;
	LAYER met2 ;
		ENCLOSURE 0.055 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
		SPACING 0.17 BY 0.17 ;

END M1M2_PR 

VIARULE M1M2_PR_R GENERATE 
	LAYER met1 ;
		ENCLOSURE 0.055 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met2 ;
		ENCLOSURE 0.085 0.055 ;
		WIDTH 0 TO 1000 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
		SPACING 0.32 BY 0.32 ;

END M1M2_PR_R 

VIARULE M1M2_PR_M GENERATE 
	LAYER met1 ;
		ENCLOSURE 0.085 0.055 ;
		WIDTH 0 TO 1000 ;
	LAYER met2 ;
		ENCLOSURE 0.055 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
		SPACING 0.17 BY 0.17 ;

END M1M2_PR_M 

VIARULE M1M2_PR_MR GENERATE 
	LAYER met1 ;
		ENCLOSURE 0.055 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met2 ;
		ENCLOSURE 0.085 0.055 ;
		WIDTH 0 TO 1000 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
		SPACING 0.17 BY 0.17 ;

END M1M2_PR_MR 

VIARULE M1M2_PR_C GENERATE 
	LAYER met1 ;
		ENCLOSURE 0.085 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met2 ;
		ENCLOSURE 0.085 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
		SPACING 0.32 BY 0.32 ;

END M1M2_PR_C 

VIARULE M2M3_PR GENERATE 
	LAYER met2 ;
		ENCLOSURE 0.04 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met3 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M2M3_PR 

VIARULE M2M3_PR_R GENERATE 
	LAYER met2 ;
		ENCLOSURE 0.085 0.04 ;
		WIDTH 0 TO 1000 ;
	LAYER met3 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M2M3_PR_R 

VIARULE M2M3_PR_M GENERATE 
	LAYER met2 ;
		ENCLOSURE 0.04 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met3 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M2M3_PR_M 

VIARULE M2M3_PR_MR GENERATE 
	LAYER met2 ;
		ENCLOSURE 0.085 0.04 ;
		WIDTH 0 TO 1000 ;
	LAYER met3 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M2M3_PR_MR 

VIARULE M2M3_PR_C GENERATE 
	LAYER met2 ;
		ENCLOSURE 0.085 0.085 ;
		WIDTH 0 TO 1000 ;
	LAYER met3 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M2M3_PR_C 

VIARULE M3M4_PR GENERATE 
	LAYER met3 ;
		ENCLOSURE 0.09 0.06 ;
		WIDTH 0 TO 1000 ;
	LAYER met4 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M3M4_PR 

VIARULE M3M4_PR_R GENERATE 
	LAYER met3 ;
		ENCLOSURE 0.06 0.09 ;
		WIDTH 0 TO 1000 ;
	LAYER met4 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M3M4_PR_R 

VIARULE M3M4_PR_M GENERATE 
	LAYER met3 ;
		ENCLOSURE 0.09 0.06 ;
		WIDTH 0 TO 1000 ;
	LAYER met4 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M3M4_PR_M 

VIARULE M3M4_PR_MR GENERATE 
	LAYER met3 ;
		ENCLOSURE 0.06 0.09 ;
		WIDTH 0 TO 1000 ;
	LAYER met4 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M3M4_PR_MR 

VIARULE M3M4_PR_C GENERATE 
	LAYER met3 ;
		ENCLOSURE 0.09 0.09 ;
		WIDTH 0 TO 1000 ;
	LAYER met4 ;
		ENCLOSURE 0.065 0.065 ;
		WIDTH 0 TO 1000 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
		SPACING 0.4 BY 0.4 ;

END M3M4_PR_C 

VIARULE M4M5_PR GENERATE 
	LAYER met4 ;
		ENCLOSURE 0.19 0.19 ;
		WIDTH 0 TO 1000 ;
	LAYER met5 ;
		ENCLOSURE 0.31 0.31 ;
		WIDTH 0 TO 1000 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
		SPACING 1.6 BY 1.6 ;

END M4M5_PR 

VIARULE M4M5_PR_R GENERATE 
	LAYER met4 ;
		ENCLOSURE 0.19 0.19 ;
		WIDTH 0 TO 1000 ;
	LAYER met5 ;
		ENCLOSURE 0.31 0.31 ;
		WIDTH 0 TO 1000 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
		SPACING 1.6 BY 1.6 ;

END M4M5_PR_R 

VIARULE M4M5_PR_M GENERATE 
	LAYER met4 ;
		ENCLOSURE 0.19 0.19 ;
		WIDTH 0 TO 1000 ;
	LAYER met5 ;
		ENCLOSURE 0.31 0.31 ;
		WIDTH 0 TO 1000 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
		SPACING 1.6 BY 1.6 ;

END M4M5_PR_M 

VIARULE M4M5_PR_MR GENERATE 
	LAYER met4 ;
		ENCLOSURE 0.19 0.19 ;
		WIDTH 0 TO 1000 ;
	LAYER met5 ;
		ENCLOSURE 0.31 0.31 ;
		WIDTH 0 TO 1000 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
		SPACING 1.6 BY 1.6 ;

END M4M5_PR_MR 

VIARULE M4M5_PR_C GENERATE 
	LAYER met4 ;
		ENCLOSURE 0.19 0.19 ;
		WIDTH 0 TO 1000 ;
	LAYER met5 ;
		ENCLOSURE 0.31 0.31 ;
		WIDTH 0 TO 1000 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
		SPACING 1.6 BY 1.6 ;

END M4M5_PR_C 

VIA M1M2_PR DEFAULT 
	RESISTANCE 4.5 ;
	LAYER met1 ;
		RECT -0.16 -0.13 0.16 0.13 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER met2 ;
		RECT -0.13 -0.16 0.13 0.16 ;

END M1M2_PR 

VIA M1M2_PR_C DEFAULT 
	RESISTANCE 4.5 ;
	LAYER met1 ;
		RECT -0.16 -0.16 0.16 0.16 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER met2 ;
		RECT -0.16 -0.16 0.16 0.16 ;

END M1M2_PR_C 

VIA M1M2_PR_M DEFAULT 
	RESISTANCE 4.5 ;
	LAYER met1 ;
		RECT -0.16 -0.13 0.16 0.13 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER met2 ;
		RECT -0.13 -0.16 0.13 0.16 ;

END M1M2_PR_M 

VIA M1M2_PR_MR DEFAULT 
	RESISTANCE 4.5 ;
	LAYER met1 ;
		RECT -0.13 -0.16 0.13 0.16 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER met2 ;
		RECT -0.13 -0.16 0.13 0.16 ;

END M1M2_PR_MR 

VIA M1M2_PR_R DEFAULT 
	RESISTANCE 4.5 ;
	LAYER met1 ;
		RECT -0.13 -0.16 0.13 0.16 ;
	LAYER via ;
		RECT -0.075 -0.075 0.075 0.075 ;
	LAYER met2 ;
		RECT -0.16 -0.13 0.16 0.13 ;

END M1M2_PR_R 

VIA M2M3_PR DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met2 ;
		RECT -0.14 -0.185 0.14 0.185 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met3 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M2M3_PR 

VIA M2M3_PR_C DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met2 ;
		RECT -0.185 -0.185 0.185 0.185 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met3 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M2M3_PR_C 

VIA M2M3_PR_M DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met2 ;
		RECT -0.14 -0.185 0.14 0.185 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met3 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M2M3_PR_M 

VIA M2M3_PR_MR DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met2 ;
		RECT -0.185 -0.14 0.185 0.14 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met3 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M2M3_PR_MR 

VIA M2M3_PR_R DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met2 ;
		RECT -0.185 -0.14 0.185 0.14 ;
	LAYER via2 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met3 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M2M3_PR_R 

VIA M3M4_PR DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met3 ;
		RECT -0.19 -0.16 0.19 0.16 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met4 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M3M4_PR 

VIA M3M4_PR_C DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met3 ;
		RECT -0.19 -0.19 0.19 0.19 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met4 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M3M4_PR_C 

VIA M3M4_PR_M DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met3 ;
		RECT -0.19 -0.16 0.19 0.16 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met4 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M3M4_PR_M 

VIA M3M4_PR_MR DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met3 ;
		RECT -0.16 -0.19 0.16 0.19 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met4 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M3M4_PR_MR 

VIA M3M4_PR_R DEFAULT 
	RESISTANCE 3.41 ;
	LAYER met3 ;
		RECT -0.16 -0.19 0.16 0.19 ;
	LAYER via3 ;
		RECT -0.1 -0.1 0.1 0.1 ;
	LAYER met4 ;
		RECT -0.165 -0.165 0.165 0.165 ;

END M3M4_PR_R 

VIA M4M5_PR DEFAULT 
	RESISTANCE 0.38 ;
	LAYER met4 ;
		RECT -0.59 -0.59 0.59 0.59 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
	LAYER met5 ;
		RECT -0.71 -0.71 0.71 0.71 ;

END M4M5_PR 

VIA M4M5_PR_C DEFAULT 
	RESISTANCE 0.38 ;
	LAYER met4 ;
		RECT -0.59 -0.59 0.59 0.59 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
	LAYER met5 ;
		RECT -0.71 -0.71 0.71 0.71 ;

END M4M5_PR_C 

VIA M4M5_PR_M DEFAULT 
	RESISTANCE 0.38 ;
	LAYER met4 ;
		RECT -0.59 -0.59 0.59 0.59 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
	LAYER met5 ;
		RECT -0.71 -0.71 0.71 0.71 ;

END M4M5_PR_M 

VIA M4M5_PR_MR DEFAULT 
	RESISTANCE 0.38 ;
	LAYER met4 ;
		RECT -0.59 -0.59 0.59 0.59 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
	LAYER met5 ;
		RECT -0.71 -0.71 0.71 0.71 ;

END M4M5_PR_MR 

VIA M4M5_PR_R DEFAULT 
	RESISTANCE 0.38 ;
	LAYER met4 ;
		RECT -0.59 -0.59 0.59 0.59 ;
	LAYER via4 ;
		RECT -0.4 -0.4 0.4 0.4 ;
	LAYER met5 ;
		RECT -0.71 -0.71 0.71 0.71 ;

END M4M5_PR_R 

SITE CoreSite 
	CLASS CORE ;
	SYMMETRY X Y ;
	SIZE 0.46 BY 4.14 ;
END CoreSite 

SITE IOSite 
	CLASS PAD ;
	SYMMETRY X Y R90 ;
	SIZE 1.0 BY 240.0 ;
END IOSite 

SITE CornerSite 
	CLASS PAD ;
	SYMMETRY X Y R90 ;
	SIZE 240.0 BY 240.0 ;
END CornerSite 

MACRO AOI221X1
	CLASS CORE ;
	FOREIGN AOI221X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.8 0.64 3.06 3.215 ;
			RECT 2.63 0.64 3.06 2.525 ;
			RECT 0.975 0.64 3.06 0.87 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.81 0.59 2.05 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.325 1.05 2.565 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.325 1.97 2.565 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.15 1.51 2.39 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.13 2.43 2.37 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.650441 LAYER met1  ;
		ANTENNAMAXAREACAR 0.552875 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 2.83 2.645 3.06 ;
			RECT 0.115 3.27 2.125 3.5 ;

	END

END AOI221X1

MACRO SDFFX1
	CLASS CORE ;
	FOREIGN SDFFX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 10.58 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.045 0.68 9.39 3.455 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.905 0.675 10.25 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.435 2.43 1.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.15 1.05 3.39 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.13968 LAYER met1  ;
		ANTENNAMAXAREACAR 1.06048 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.82 2.43 3.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 10.58 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 10.58 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.675 3.375 5.715 3.605 ;
			RECT 5.485 2.475 5.715 3.605 ;
			RECT 3.675 0.705 3.905 3.605 ;
			RECT 1.435 3.375 3.475 3.605 ;
			RECT 3.245 0.705 3.475 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 8.585 0.88 8.815 3.53 ;
			RECT 7.725 0.68 7.955 3.53 ;
			RECT 6.775 1.145 7.005 2.795 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.915 0.705 6.145 3.235 ;
			RECT 4.965 0.705 5.195 3.235 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFX1

MACRO OR3X2
	CLASS CORE ;
	FOREIGN OR3X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.925 3.24 2.43 3.53 ;
			RECT 2.17 0.535 2.43 3.53 ;
			RECT 1.925 0.535 2.43 0.825 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.46 1.51 2.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.06 1.05 2.3 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.742857 LAYER met1  ;
		ANTENNAMAXAREACAR 0.631429 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.31 0.59 2.55 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.87 1.2 3.5 ;
			RECT 0.97 2.87 2.03 3.1 ;
			RECT 1.8 1.09 2.03 3.1 ;
			RECT 1.36 1.09 2.03 1.32 ;
			RECT 1.36 0.475 1.59 1.32 ;
			RECT 0.115 0.475 1.59 0.705 ;

	END

END OR3X2

MACRO OAI211X1
	CLASS CORE ;
	FOREIGN OAI211X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.99 2.865 2.43 3.125 ;
			RECT 2.17 0.61 2.43 3.125 ;
			RECT 1.85 0.61 2.43 0.905 ;
			RECT 1.865 2.865 2.095 3.53 ;
			RECT 0.99 2.865 1.25 3.515 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.19 0.59 2.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.285 1.05 2.525 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.402116 LAYER met1  ;
		ANTENNAMAXAREACAR 0.341799 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.31 1.51 2.55 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.42328 LAYER met1  ;
		ANTENNAMAXAREACAR 0.359788 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.32 1.97 2.56 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.419753 LAYER met1  ;
		ANTENNAMAXAREACAR 0.35679 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.005 0.61 1.235 0.935 ;
			RECT 0.145 0.61 0.375 0.935 ;
			RECT 0.145 0.61 1.235 0.84 ;

	END

END OAI211X1

MACRO AOI222X1
	CLASS CORE ;
	FOREIGN AOI222X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.14 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.245 0.68 3.475 1.33 ;
			RECT 0.975 0.68 3.475 0.91 ;
			RECT 2.63 0.68 3.045 3.09 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.05 0.59 2.29 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.444444 LAYER met1  ;
		ANTENNAMAXAREACAR 0.377778 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.495 1.05 2.735 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.444444 LAYER met1  ;
		ANTENNAMAXAREACAR 0.377778 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.49 1.97 2.73 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.567901 LAYER met1  ;
		ANTENNAMAXAREACAR 0.482716 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.1 1.51 2.34 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.444444 LAYER met1  ;
		ANTENNAMAXAREACAR 0.377778 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.33 2.43 2.57 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.617284 LAYER met1  ;
		ANTENNAMAXAREACAR 0.524691 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.765 3.81 3.005 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.70194 LAYER met1  ;
		ANTENNAMAXAREACAR 0.596649 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.14 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.14 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 3.27 3.505 3.5 ;
			RECT 0.115 2.9 2.125 3.13 ;

	END

END AOI222X1

MACRO AND4X2
	CLASS CORE ;
	FOREIGN AND4X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.355 3.24 2.89 3.53 ;
			RECT 2.63 0.61 2.89 3.53 ;
			RECT 2.355 0.61 2.89 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.425 1.97 2.665 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.02222 LAYER met1  ;
		ANTENNAMAXAREACAR 0.868889 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.865 1.51 3.105 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.968889 LAYER met1  ;
		ANTENNAMAXAREACAR 0.823556 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.055 1.05 2.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.920635 LAYER met1  ;
		ANTENNAMAXAREACAR 0.78254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.055 0.59 2.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.920635 LAYER met1  ;
		ANTENNAMAXAREACAR 0.78254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.545 3.27 2.125 3.5 ;
			RECT 1.895 2.87 2.125 3.5 ;
			RECT 1.895 2.87 2.48 3.1 ;
			RECT 2.215 1.04 2.445 3.1 ;
			RECT 2.21 2.0 2.445 2.29 ;
			RECT 1.985 0.64 2.215 1.27 ;
			RECT 0.115 0.64 2.215 0.87 ;

	END

END AND4X2

MACRO AND2X2
	CLASS CORE ;
	FOREIGN AND2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.495 3.18 1.97 3.47 ;
			RECT 1.71 0.655 1.97 3.47 ;
			RECT 1.495 0.655 1.97 0.945 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 0.0007 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.00023 LAYER met1  ;
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.535 1.51 2.775 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.26222 LAYER met1  ;
		ANTENNAMAXAREACAR 1.07289 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.745 0.59 2.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.910476 LAYER met1  ;
		ANTENNAMAXAREACAR 0.773905 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 3.24 0.99 3.53 ;
			RECT 0.76 0.685 0.99 3.53 ;
			RECT 0.145 0.655 0.375 0.945 ;
			RECT 0.145 0.685 0.99 0.915 ;

	END

END AND2X2

MACRO NOR3X4
	CLASS CORE ;
	FOREIGN NOR3X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.44 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.105 3.27 6.11 3.5 ;
			RECT 5.825 0.61 6.11 3.5 ;
			RECT 0.575 0.61 6.11 0.9 ;
			RECT 4.965 2.85 5.195 3.5 ;
			RECT 4.105 2.85 4.335 3.5 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.085 1.05 2.325 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.175 1.04 2.435 2.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.258377 LAYER met1  ;
		ANTENNAMAXAREACAR 0.270591 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.04 5.19 2.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.44 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.44 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.395 2.47 5.625 3.12 ;
			RECT 4.535 2.47 4.765 3.12 ;
			RECT 3.155 2.47 3.385 3.12 ;
			RECT 2.295 2.47 2.525 3.12 ;
			RECT 2.295 2.47 5.625 2.7 ;
			RECT 0.145 3.27 3.815 3.5 ;
			RECT 3.585 2.85 3.815 3.5 ;
			RECT 2.725 2.85 2.955 3.5 ;
			RECT 1.865 2.49 2.095 3.5 ;
			RECT 1.005 2.49 1.235 3.5 ;
			RECT 0.145 2.49 0.375 3.5 ;

	END

END NOR3X4

MACRO DFFRX1
	CLASS CORE ;
	FOREIGN DFFRX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 9.2 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 7.69 2.44 7.955 3.45 ;
			RECT 7.69 0.68 7.955 1.33 ;
			RECT 7.69 0.68 7.95 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 8.585 2.44 8.87 3.45 ;
			RECT 8.61 0.68 8.87 3.45 ;
			RECT 8.585 0.68 8.87 1.33 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.315 1.05 3.555 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.07937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.91746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.385 1.05 1.625 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 6.77 1.405 7.03 2.645 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.9746 LAYER met1  ;
		ANTENNAMAXAREACAR 2.62016 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END RN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 9.2 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 9.2 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 6.345 0.765 6.575 3.53 ;
			RECT 5.915 0.765 6.575 0.995 ;
			RECT 5.915 0.705 6.145 0.995 ;
			RECT 1.435 3.375 3.905 3.605 ;
			RECT 3.675 2.505 3.905 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 2.725 2.945 2.955 3.235 ;
			RECT 1.865 2.945 2.095 3.235 ;
			RECT 1.865 3.005 2.955 3.175 ;
			RECT 7.205 0.61 7.435 3.53 ;
			RECT 4.965 1.145 5.195 2.795 ;
			RECT 4.535 0.705 4.765 3.235 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 3.245 0.705 3.475 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFRX1

MACRO SDFFRX1
	CLASS CORE ;
	FOREIGN SDFFRX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 11.5 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.825 0.685 11.17 3.455 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.965 0.68 10.25 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.4 2.43 1.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.125 1.05 3.365 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.660317 LAYER met1  ;
		ANTENNAMAXAREACAR 0.56127 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.17 5.19 2.41 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.28571 LAYER met1  ;
		ANTENNAMAXAREACAR 2.0346 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END RN
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.16508 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08206 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.78 2.43 3.02 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 11.5 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 11.5 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 9.45 0.765 9.68 3.235 ;
			RECT 8.985 0.765 9.68 0.935 ;
			RECT 8.585 0.705 8.815 3.235 ;
			RECT 8.495 0.705 8.815 0.995 ;
			RECT 6.775 0.705 7.005 3.235 ;
			RECT 6.775 1.855 7.545 2.085 ;
			RECT 3.675 3.375 6.145 3.605 ;
			RECT 5.915 2.475 6.145 3.605 ;
			RECT 3.675 0.705 3.905 3.605 ;
			RECT 1.435 3.57 3.475 3.8 ;
			RECT 3.245 0.705 3.475 3.8 ;
			RECT 1.435 0.705 1.665 3.8 ;
			RECT 0.15 0.71 0.38 3.24 ;
			RECT 0.145 2.945 0.38 3.235 ;
			RECT 0.145 2.505 0.38 2.795 ;
			RECT 0.145 1.145 0.38 1.435 ;
			RECT 0.145 0.705 0.375 0.995 ;
			RECT 7.715 1.145 7.945 2.795 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.485 0.705 5.715 3.235 ;
			RECT 4.075 3.005 5.225 3.175 ;
			RECT 2.725 0.705 2.955 3.235 ;

	END

END SDFFRX1

MACRO OAI22X2
	CLASS CORE ;
	FOREIGN OAI22X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.105 0.87 4.335 3.45 ;
			RECT 2.385 2.71 4.335 2.94 ;
			RECT 4.01 0.87 4.335 2.94 ;
			RECT 3.675 0.87 4.335 1.16 ;
			RECT 1.435 0.87 4.335 1.1 ;
			RECT 3.245 2.71 3.475 3.0 ;
			RECT 2.385 2.71 2.615 3.0 ;
			RECT 1.435 0.87 1.665 1.16 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.545 0.59 2.785 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.24 2.89 2.48 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.585 1.51 2.825 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.333333 LAYER met1  ;
		ANTENNAMAXAREACAR 0.361111 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.325 3.81 2.565 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.005 0.44 1.235 1.09 ;
			RECT 0.145 0.44 0.375 1.09 ;
			RECT 4.105 0.44 4.335 0.73 ;
			RECT 3.245 0.44 3.475 0.73 ;
			RECT 2.385 0.44 2.615 0.73 ;
			RECT 1.865 0.44 2.095 0.73 ;
			RECT 0.145 0.44 4.335 0.67 ;
			RECT 3.675 3.14 3.905 3.43 ;
			RECT 1.435 3.14 3.905 3.37 ;
			RECT 1.435 3.08 1.665 3.37 ;
			RECT 0.575 3.57 3.045 3.8 ;
			RECT 2.815 3.51 3.045 3.8 ;
			RECT 0.575 3.51 0.805 3.8 ;

	END

END OAI22X2

MACRO DFFX4
	CLASS CORE ;
	FOREIGN DFFX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 10.58 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 8.125 0.68 8.45 3.45 ;
			RECT 7.265 1.77 8.45 2.0 ;
			RECT 7.265 0.68 7.495 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.845 0.68 10.25 3.45 ;
			RECT 8.985 1.77 10.25 2.0 ;
			RECT 8.985 0.68 9.215 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.655 1.05 1.895 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 10.58 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 10.58 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.485 3.42 3.715 ;
			RECT 3.19 0.415 3.42 3.715 ;
			RECT 1.435 2.945 1.665 3.715 ;
			RECT 1.435 0.415 1.665 0.995 ;
			RECT 1.435 0.415 3.42 0.645 ;
			RECT 6.405 0.68 6.635 3.45 ;
			RECT 5.455 0.745 5.685 3.315 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 2.725 0.785 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFX4

MACRO XNOR2X2
	CLASS CORE ;
	FOREIGN XNOR2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 2.44 3.015 3.09 ;
			RECT 2.63 0.61 3.015 1.26 ;
			RECT 2.63 0.61 2.89 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.175 1.05 2.415 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.679365 LAYER met1  ;
		ANTENNAMAXAREACAR 0.57746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.09 0.59 2.33 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.930159 LAYER met1  ;
		ANTENNAMAXAREACAR 0.882381 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.3 3.415 3.47 ;
			RECT 3.245 1.65 3.415 3.47 ;
			RECT 1.435 3.18 1.795 3.47 ;
			RECT 1.655 0.44 1.795 3.47 ;
			RECT 3.215 1.65 3.445 1.94 ;
			RECT 1.435 0.44 1.795 0.73 ;
			RECT 1.935 2.505 2.165 2.795 ;
			RECT 2.025 1.225 2.165 2.795 ;
			RECT 1.935 1.225 2.165 1.515 ;
			RECT 1.005 3.18 1.235 3.47 ;
			RECT 1.05 2.8 1.19 3.47 ;
			RECT 1.05 2.8 1.475 2.94 ;
			RECT 1.335 0.895 1.475 2.94 ;
			RECT 1.19 1.655 1.475 1.945 ;
			RECT 1.05 0.895 1.475 1.035 ;
			RECT 1.05 0.44 1.19 1.035 ;
			RECT 1.005 0.44 1.235 0.73 ;
			RECT 0.01 3.45 0.375 3.74 ;
			RECT 0.01 0.425 0.18 3.74 ;
			RECT 0.01 2.505 0.29 2.795 ;
			RECT 0.01 0.425 0.375 0.715 ;

	END

END XNOR2X2

MACRO INVX2
	CLASS CORE ;
	FOREIGN INVX2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 2.735 1.05 3.385 ;
			RECT 0.79 0.61 1.05 3.385 ;
			RECT 0.575 0.61 1.05 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.29 0.59 2.53 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.382716 LAYER met1  ;
		ANTENNAMAXAREACAR 0.376279 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD

END INVX2

MACRO BUFX4
	CLASS CORE ;
	FOREIGN BUFX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.005 3.24 2.095 3.53 ;
			RECT 1.71 2.88 2.095 3.53 ;
			RECT 1.71 0.61 2.095 1.26 ;
			RECT 1.71 0.61 1.97 3.53 ;
			RECT 1.005 0.615 2.095 0.905 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.165 1.05 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.723104 LAYER met1  ;
		ANTENNAMAXAREACAR 0.614638 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 1.04 0.375 2.73 ;

	END

END BUFX4

MACRO XOR2X1
	CLASS CORE ;
	FOREIGN XOR2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.785 2.48 3.35 2.74 ;
			RECT 3.09 1.005 3.35 2.74 ;
			RECT 2.77 1.005 3.35 1.265 ;
			RECT 2.77 0.615 3.03 1.265 ;
			RECT 2.785 2.48 3.015 3.49 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.48 1.05 2.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.819048 LAYER met1  ;
		ANTENNAMAXAREACAR 0.69619 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 2.05 0.59 3.29 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.00952 LAYER met1  ;
		ANTENNAMAXAREACAR 1.97794 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 3.32 2.57 3.49 ;
			RECT 2.31 0.575 2.57 3.49 ;
			RECT 1.405 0.535 2.565 0.705 ;
			RECT 0.975 2.98 2.075 3.15 ;
			RECT 1.815 0.845 2.075 3.15 ;
			RECT 0.975 0.845 2.075 1.015 ;
			RECT 0.01 3.435 0.375 3.725 ;
			RECT 0.01 0.655 0.18 3.725 ;
			RECT 0.01 1.61 0.29 1.9 ;
			RECT 0.01 0.655 0.375 0.945 ;

	END

END XOR2X1

MACRO NOR4X1
	CLASS CORE ;
	FOREIGN NOR4X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.865 3.235 2.43 3.525 ;
			RECT 2.17 0.625 2.43 3.525 ;
			RECT 0.145 0.625 2.43 0.915 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 0.0014 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.00046 LAYER met1  ;
	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.685 0.59 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.165 1.05 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.514991 LAYER met1  ;
		ANTENNAMAXAREACAR 0.437743 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.685 1.51 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.536155 LAYER met1  ;
		ANTENNAMAXAREACAR 0.455732 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.205 1.97 2.445 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.557319 LAYER met1  ;
		ANTENNAMAXAREACAR 0.473721 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD

END NOR4X1

MACRO NOR2X1
	CLASS CORE ;
	FOREIGN NOR2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.84 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.105 2.5 1.51 3.51 ;
			RECT 1.25 0.62 1.51 3.51 ;
			RECT 0.635 0.62 1.51 0.91 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.76 0.59 3.0 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.391534 LAYER met1  ;
		ANTENNAMAXAREACAR 0.332804 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.125 1.05 2.365 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.405644 LAYER met1  ;
		ANTENNAMAXAREACAR 0.344797 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.84 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.84 4.34 ;

		END 

	END VDD

END NOR2X1

MACRO NAND3X2
	CLASS CORE ;
	FOREIGN NAND3X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.545 3.27 3.045 3.5 ;
			RECT 2.63 2.49 3.045 3.5 ;
			RECT 2.63 1.025 3.045 1.315 ;
			RECT 2.63 1.025 2.89 3.5 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.65 0.59 2.89 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.405644 LAYER met1  ;
		ANTENNAMAXAREACAR 0.395767 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.65 1.51 2.89 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.38448 LAYER met1  ;
		ANTENNAMAXAREACAR 0.377778 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.53 2.43 2.77 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.442681 LAYER met1  ;
		ANTENNAMAXAREACAR 0.427249 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 0.64 3.505 0.87 ;
			RECT 0.115 1.025 2.125 1.255 ;

	END

END NAND3X2

MACRO DFFSX4
	CLASS CORE ;
	FOREIGN DFFSX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 11.96 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.445 0.68 9.79 3.45 ;
			RECT 8.585 1.77 9.79 2.0 ;
			RECT 8.585 0.68 8.815 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.885 2.44 11.395 3.45 ;
			RECT 10.885 0.68 11.395 1.33 ;
			RECT 10.885 0.68 11.17 3.45 ;
			RECT 10.305 1.77 11.17 2.0 ;
			RECT 10.305 0.68 10.535 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.655 1.05 1.895 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.5 3.35 2.74 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.94286 LAYER met1  ;
		ANTENNAMAXAREACAR 1.74318 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 11.96 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 11.96 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.825 2.945 6.055 3.235 ;
			RECT 4.965 2.945 5.195 3.235 ;
			RECT 4.965 3.005 6.055 3.175 ;
			RECT 3.215 3.355 4.335 3.585 ;
			RECT 4.105 0.705 4.335 3.585 ;
			RECT 2.295 0.705 2.525 1.795 ;
			RECT 2.295 0.705 4.335 0.935 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 1.435 2.965 3.905 3.195 ;
			RECT 3.675 2.505 3.905 3.195 ;
			RECT 7.725 0.68 7.955 3.45 ;
			RECT 6.775 0.745 7.005 3.315 ;
			RECT 4.965 1.145 5.195 2.795 ;
			RECT 4.535 0.705 4.765 3.235 ;
			RECT 2.71 1.145 2.94 2.795 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFSX4

MACRO SDFFSX4
	CLASS CORE ;
	FOREIGN SDFFSX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 14.26 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 11.685 0.68 12.09 3.45 ;
			RECT 10.825 1.77 12.09 2.0 ;
			RECT 10.825 0.68 11.055 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 13.405 0.675 13.93 3.45 ;
			RECT 12.545 1.77 13.93 2.0 ;
			RECT 12.545 0.68 12.775 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.435 2.43 1.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.15 1.05 3.39 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.16508 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08206 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.82 2.43 3.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.39 1.485 5.65 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.90794 LAYER met1  ;
		ANTENNAMAXAREACAR 1.71349 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 14.265 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 14.265 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.485 3.005 6.575 3.235 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.485 2.945 5.715 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 5.915 0.705 6.145 2.795 ;
			RECT 3.675 0.705 6.145 0.935 ;
			RECT 1.435 3.375 3.475 3.605 ;
			RECT 3.245 0.705 3.475 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 9.965 0.68 10.195 3.45 ;
			RECT 9.015 0.88 9.245 3.315 ;
			RECT 7.175 2.975 8.325 3.205 ;
			RECT 7.205 1.145 7.435 2.795 ;
			RECT 6.775 0.705 7.005 3.235 ;
			RECT 4.965 1.145 5.195 3.235 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFSX4

MACRO CLKINVX2
	CLASS CORE ;
	FOREIGN CLKINVX2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.235 1.05 3.525 ;
			RECT 0.79 0.61 1.05 3.525 ;
			RECT 0.575 0.61 1.05 1.26 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.54 0.59 2.78 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.326279 LAYER met1  ;
		ANTENNAMAXAREACAR 0.328307 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD

END CLKINVX2

MACRO OAI21X2
	CLASS CORE ;
	FOREIGN OAI21X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.245 2.73 3.475 3.38 ;
			RECT 3.09 1.1 3.35 3.1 ;
			RECT 1.435 2.87 3.475 3.1 ;
			RECT 1.435 1.1 3.35 1.33 ;
			RECT 2.385 2.87 2.615 3.365 ;
			RECT 1.435 2.87 1.665 3.365 ;
			RECT 1.435 1.04 1.665 1.33 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.055 0.59 2.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.47 2.89 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.47 1.51 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.245 0.61 3.475 0.9 ;
			RECT 2.385 0.61 2.615 0.9 ;
			RECT 1.865 0.61 2.095 0.9 ;
			RECT 1.005 0.61 1.235 0.9 ;
			RECT 0.145 0.61 0.375 0.9 ;
			RECT 0.145 0.61 3.475 0.84 ;
			RECT 0.575 3.52 3.045 3.75 ;
			RECT 2.815 3.24 3.045 3.75 ;
			RECT 0.575 2.52 0.805 3.75 ;

	END

END OAI21X2

MACRO CLKBUFX4
	CLASS CORE ;
	FOREIGN CLKBUFX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.005 3.225 2.43 3.515 ;
			RECT 2.17 0.61 2.43 3.515 ;
			RECT 1.865 2.505 2.43 3.515 ;
			RECT 1.865 0.61 2.43 1.26 ;
			RECT 1.005 0.61 2.43 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.635 1.05 2.875 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.666667 LAYER met1  ;
		ANTENNAMAXAREACAR 0.566667 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 0.61 0.375 3.515 ;
			RECT 1.26 1.11 1.52 1.77 ;
			RECT 0.145 1.11 1.52 1.37 ;

	END

END CLKBUFX4

MACRO XOR2X4
	CLASS CORE ;
	FOREIGN XOR2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.52 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.655 2.465 5.19 2.755 ;
			RECT 4.93 0.695 5.19 2.755 ;
			RECT 3.795 1.77 5.19 2.0 ;
			RECT 4.655 0.695 5.19 0.985 ;
			RECT 3.795 0.68 4.025 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 2.09 0.59 3.33 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.07 1.05 2.31 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.478458 LAYER met1  ;
		ANTENNAMAXAREACAR 0.472222 LAYER met1  ;
		ANTENNAGATEAREA 0.441 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.52 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.52 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.985 1.32 2.215 3.09 ;
			RECT 1.985 1.51 3.595 1.74 ;
			RECT 1.615 1.01 1.845 2.29 ;
			RECT 1.615 1.01 2.675 1.18 ;
			RECT 1.005 2.945 1.36 3.235 ;
			RECT 1.19 0.46 1.36 3.235 ;
			RECT 1.19 1.66 1.42 1.95 ;
			RECT 1.005 0.46 1.36 0.75 ;
			RECT 0.01 3.475 0.375 3.765 ;
			RECT 0.01 0.46 0.18 3.765 ;
			RECT 0.01 1.66 0.24 1.95 ;
			RECT 0.01 0.46 0.375 0.75 ;
			RECT 1.525 0.64 3.195 0.87 ;

	END

END XOR2X4

MACRO AND3X2
	CLASS CORE ;
	FOREIGN AND3X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.925 3.095 2.43 3.385 ;
			RECT 2.17 0.61 2.43 3.385 ;
			RECT 1.925 0.61 2.43 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.105 1.51 2.345 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.692063 LAYER met1  ;
		ANTENNAMAXAREACAR 0.588254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.44 1.05 1.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.634921 LAYER met1  ;
		ANTENNAMAXAREACAR 0.539683 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.945 1.05 3.185 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.23048 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0459 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 3.36 1.285 3.53 ;
			RECT 0.145 0.705 0.375 3.53 ;

	END

END AND3X2

MACRO NOR4X4
	CLASS CORE ;
	FOREIGN NOR4X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.82 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 0.61 7.82 0.9 ;
			RECT 7.23 0.61 7.49 2.97 ;
			RECT 7.1 2.71 7.36 3.36 ;
			RECT 6.255 0.61 6.485 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.045 1.05 2.285 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.175 1.05 2.435 2.29 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.258377 LAYER met1  ;
		ANTENNAMAXAREACAR 0.270591 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 1.065 4.73 2.305 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.248677 LAYER met1  ;
		ANTENNAMAXAREACAR 0.262346 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 6.77 1.105 7.03 2.345 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.82 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.82 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.105 3.5 7.775 3.73 ;
			RECT 7.545 3.24 7.775 3.73 ;
			RECT 6.685 2.49 6.915 3.73 ;
			RECT 5.825 2.49 6.055 3.73 ;
			RECT 4.965 2.85 5.195 3.73 ;
			RECT 4.105 2.85 4.335 3.73 ;
			RECT 5.395 2.47 5.625 3.12 ;
			RECT 4.535 2.47 4.765 3.12 ;
			RECT 3.155 2.47 3.385 3.12 ;
			RECT 2.295 2.47 2.525 3.12 ;
			RECT 2.295 2.47 5.625 2.7 ;
			RECT 0.145 3.27 3.815 3.5 ;
			RECT 3.585 2.85 3.815 3.5 ;
			RECT 2.725 2.85 2.955 3.5 ;
			RECT 1.865 2.49 2.095 3.5 ;
			RECT 1.005 2.49 1.235 3.5 ;
			RECT 0.145 2.49 0.375 3.5 ;

	END

END NOR4X4

MACRO NOR2X4
	CLASS CORE ;
	FOREIGN NOR2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.14 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.155 2.44 3.385 3.09 ;
			RECT 0.575 0.61 3.385 0.9 ;
			RECT 2.17 2.44 3.385 2.67 ;
			RECT 2.17 0.61 2.525 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.405 0.59 2.645 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.314815 LAYER met1  ;
		ANTENNAMAXAREACAR 0.344048 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.555 3.81 2.795 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.346561 LAYER met1  ;
		ANTENNAMAXAREACAR 0.371032 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.14 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.14 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 3.845 3.5 ;

	END

END NOR2X4

MACRO DFFSX1
	CLASS CORE ;
	FOREIGN DFFSX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 9.2 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 7.69 2.44 7.955 3.45 ;
			RECT 7.69 0.68 7.955 1.33 ;
			RECT 7.69 0.68 7.95 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 8.585 0.68 8.87 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.655 1.05 1.895 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 3.085 1.5 3.345 2.74 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.94603 LAYER met1  ;
		ANTENNAMAXAREACAR 1.74587 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 9.2 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 9.2 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.825 2.945 6.055 3.235 ;
			RECT 4.965 2.945 5.195 3.235 ;
			RECT 4.965 2.945 6.055 3.175 ;
			RECT 3.215 3.355 4.335 3.585 ;
			RECT 4.105 0.705 4.335 3.585 ;
			RECT 2.295 0.705 2.525 1.795 ;
			RECT 2.295 0.705 4.335 0.935 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 1.435 2.965 3.905 3.195 ;
			RECT 3.675 2.505 3.905 3.195 ;
			RECT 7.205 0.705 7.435 3.235 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 4.965 1.145 5.195 2.795 ;
			RECT 4.535 0.705 4.765 3.235 ;
			RECT 2.685 1.145 2.915 2.795 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFSX1

MACRO SDFFSX1
	CLASS CORE ;
	FOREIGN SDFFSX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 11.5 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.965 0.68 10.31 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.825 0.675 11.17 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.435 2.43 1.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.15 1.05 3.39 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.16508 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08206 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.82 2.43 3.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.39 1.485 5.65 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.90794 LAYER met1  ;
		ANTENNAMAXAREACAR 1.71349 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 11.5 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 11.5 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.485 3.005 6.575 3.235 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.485 2.945 5.715 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 5.915 0.705 6.145 2.795 ;
			RECT 3.675 0.705 6.145 0.935 ;
			RECT 1.435 3.375 3.475 3.605 ;
			RECT 3.245 0.705 3.475 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 9.445 0.705 9.675 3.235 ;
			RECT 8.585 0.705 8.815 3.235 ;
			RECT 7.175 2.975 8.325 3.205 ;
			RECT 7.205 1.145 7.435 2.795 ;
			RECT 6.775 0.705 7.005 3.235 ;
			RECT 4.965 1.145 5.195 3.235 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFSX1

MACRO DFFX1
	CLASS CORE ;
	FOREIGN DFFX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 8.28 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 6.77 0.68 7.095 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 7.69 2.44 7.955 3.45 ;
			RECT 7.69 0.68 7.955 1.33 ;
			RECT 7.69 0.68 7.95 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.655 1.05 1.895 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 8.28 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 8.28 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.485 3.42 3.715 ;
			RECT 3.19 0.415 3.42 3.715 ;
			RECT 1.435 2.945 1.665 3.715 ;
			RECT 1.435 0.415 1.665 0.995 ;
			RECT 1.435 0.415 3.42 0.645 ;
			RECT 6.345 0.68 6.575 3.45 ;
			RECT 5.395 0.745 5.625 3.315 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 2.725 0.785 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFX1

MACRO BUFX16
	CLASS CORE ;
	FOREIGN BUFX16 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 9.2 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 8.15 2.48 8.545 3.49 ;
			RECT 2.295 2.105 8.545 2.335 ;
			RECT 8.15 0.645 8.545 1.295 ;
			RECT 8.15 0.645 8.41 3.49 ;
			RECT 7.455 0.645 7.685 3.49 ;
			RECT 6.595 0.645 6.825 3.49 ;
			RECT 5.735 0.645 5.965 3.49 ;
			RECT 4.875 0.645 5.105 3.49 ;
			RECT 4.015 0.645 4.245 3.49 ;
			RECT 3.155 0.645 3.385 3.49 ;
			RECT 2.295 0.645 2.525 3.49 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.435 1.05 2.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 9.2 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 9.2 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.42 3.2 0.805 3.49 ;
			RECT 0.42 0.645 0.65 3.49 ;
			RECT 0.42 0.645 0.805 1.295 ;
			RECT 1.435 0.645 1.665 3.49 ;

	END

END BUFX16

MACRO OR4X2
	CLASS CORE ;
	FOREIGN OR4X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.355 3.24 2.89 3.53 ;
			RECT 2.63 0.535 2.89 3.53 ;
			RECT 2.355 0.535 2.89 0.825 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.47 1.97 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.768254 LAYER met1  ;
		ANTENNAMAXAREACAR 0.653016 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.145 1.51 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.72381 LAYER met1  ;
		ANTENNAMAXAREACAR 0.615238 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.435 1.05 2.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.685714 LAYER met1  ;
		ANTENNAMAXAREACAR 0.582857 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.32 1.145 0.58 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.679365 LAYER met1  ;
		ANTENNAMAXAREACAR 0.57746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.87 1.2 3.5 ;
			RECT 0.97 2.87 2.37 3.1 ;
			RECT 2.14 1.07 2.37 3.1 ;
			RECT 1.82 1.07 2.37 1.3 ;
			RECT 1.82 0.475 2.05 1.3 ;
			RECT 0.545 0.475 2.05 0.705 ;

	END

END OR4X2

MACRO OR2X2
	CLASS CORE ;
	FOREIGN OR2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.495 3.24 1.97 3.53 ;
			RECT 1.71 0.535 1.97 3.53 ;
			RECT 1.495 0.535 1.97 0.825 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.455 1.05 2.695 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.704762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.599048 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.05 0.59 2.29 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.704762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.599048 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.84 1.2 3.5 ;
			RECT 1.19 0.965 1.42 3.07 ;
			RECT 0.765 0.965 1.42 1.195 ;
			RECT 0.765 0.475 0.995 1.195 ;
			RECT 0.545 0.475 0.995 0.705 ;

	END

END OR2X2

MACRO INVX16
	CLASS CORE ;
	FOREIGN INVX16 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.36 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.545 3.21 6.855 3.5 ;
			RECT 0.545 0.61 6.855 0.9 ;
			RECT 4.01 0.61 4.27 3.5 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.465 0.59 2.705 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.307099 LAYER met1  ;
		ANTENNAMAXAREACAR 0.356603 LAYER met1  ;
		ANTENNAGATEAREA 4.536 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.36 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.36 4.34 ;

		END 

	END VDD

END INVX16

MACRO OAI222X2
	CLASS CORE ;
	FOREIGN OAI222X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.9 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.915 2.93 6.145 3.22 ;
			RECT 5.055 1.07 6.145 1.21 ;
			RECT 5.915 0.92 6.145 1.21 ;
			RECT 1.435 2.93 6.145 3.07 ;
			RECT 5.39 1.07 5.65 3.07 ;
			RECT 5.055 0.92 5.285 1.21 ;
			RECT 3.675 2.93 3.905 3.22 ;
			RECT 1.435 2.93 1.665 3.22 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.42 0.59 2.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.333333 LAYER met1  ;
		ANTENNAMAXAREACAR 0.334303 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.425 1.51 2.665 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.41 2.89 2.65 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.44 3.81 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.485 5.19 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.85 1.44 6.11 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.9 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.9 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 6.345 0.61 6.575 0.9 ;
			RECT 5.485 0.61 5.715 0.9 ;
			RECT 4.625 0.61 4.855 0.9 ;
			RECT 3.675 0.61 3.905 0.9 ;
			RECT 2.815 0.61 3.045 0.9 ;
			RECT 2.815 0.61 6.575 0.75 ;
			RECT 4.625 3.39 6.575 3.53 ;
			RECT 6.345 3.24 6.575 3.53 ;
			RECT 5.485 3.24 5.715 3.53 ;
			RECT 4.625 3.24 4.855 3.53 ;
			RECT 0.145 1.07 4.335 1.21 ;
			RECT 4.105 0.92 4.335 1.21 ;
			RECT 3.245 0.92 3.475 1.21 ;
			RECT 2.385 0.92 2.615 1.21 ;
			RECT 1.865 0.92 2.095 1.21 ;
			RECT 1.005 0.92 1.235 1.21 ;
			RECT 0.145 0.92 0.375 1.21 ;
			RECT 2.385 3.39 4.335 3.53 ;
			RECT 4.105 3.24 4.335 3.53 ;
			RECT 3.245 3.24 3.475 3.53 ;
			RECT 2.385 3.24 2.615 3.53 ;
			RECT 0.145 3.39 2.095 3.53 ;
			RECT 1.865 3.24 2.095 3.53 ;
			RECT 1.005 3.24 1.235 3.53 ;
			RECT 0.145 3.24 0.375 3.53 ;

	END

END OAI222X2

MACRO CLKMX2X2
	CLASS CORE ;
	FOREIGN CLKMX2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 0.68 3.015 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.02 1.05 3.26 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.505 2.43 2.745 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN S0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.69 1.51 2.93 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.09524 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08746 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END S0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.24 1.88 3.53 ;
			RECT 1.65 0.705 1.88 3.53 ;
			RECT 1.435 0.705 1.88 0.995 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END CLKMX2X2

MACRO NOR3X1
	CLASS CORE ;
	FOREIGN NOR3X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.435 2.865 1.97 3.155 ;
			RECT 1.71 0.61 1.97 3.155 ;
			RECT 0.575 0.61 1.97 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.165 0.59 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.685 1.05 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.514991 LAYER met1  ;
		ANTENNAMAXAREACAR 0.437743 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.4 1.51 2.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.536155 LAYER met1  ;
		ANTENNAMAXAREACAR 0.455732 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD

END NOR3X1

MACRO NAND4X2
	CLASS CORE ;
	FOREIGN NAND4X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.545 3.24 3.905 3.53 ;
			RECT 3.55 1.04 3.905 1.33 ;
			RECT 3.55 1.04 3.81 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.205 0.59 2.445 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.385 1.415 1.645 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.47 2.89 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.47 4.27 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.393298 LAYER met1  ;
		ANTENNAMAXAREACAR 0.334303 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.105 0.535 4.335 0.9 ;
			RECT 3.245 0.535 3.475 0.9 ;
			RECT 2.385 0.535 2.615 0.9 ;
			RECT 2.385 0.535 4.335 0.765 ;
			RECT 1.405 1.04 3.075 1.27 ;
			RECT 0.115 0.64 2.125 0.87 ;

	END

END NAND4X2

MACRO NAND2X2
	CLASS CORE ;
	FOREIGN NAND2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.18 1.665 3.47 ;
			RECT 1.25 2.46 1.665 3.47 ;
			RECT 1.25 1.04 1.665 1.33 ;
			RECT 1.25 1.04 1.51 3.47 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.29 0.59 2.53 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.375661 LAYER met1  ;
		ANTENNAMAXAREACAR 0.370282 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.76 1.05 3.0 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.460317 LAYER met1  ;
		ANTENNAMAXAREACAR 0.44224 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 0.59 2.125 0.76 ;

	END

END NAND2X2

MACRO DFFRX4
	CLASS CORE ;
	FOREIGN DFFRX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 12.42 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 9.875 2.44 10.25 3.45 ;
			RECT 9.99 0.68 10.25 3.45 ;
			RECT 9.015 1.77 10.25 2.0 ;
			RECT 9.875 0.68 10.25 1.33 ;
			RECT 9.015 0.68 9.245 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 11.595 2.44 12.09 3.45 ;
			RECT 11.83 0.68 12.09 3.45 ;
			RECT 10.735 1.77 12.09 2.0 ;
			RECT 11.595 0.68 12.09 1.33 ;
			RECT 10.735 0.68 10.965 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.045 1.05 3.285 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.1873 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00921 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.645 1.05 1.885 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.85 1.85 6.11 3.09 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.45156 LAYER met1  ;
		ANTENNAMAXAREACAR 1.36986 LAYER met1  ;
		ANTENNAGATEAREA 0.609 LAYER met1  ;
	END RN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 12.425 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 12.425 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 7.635 0.43 7.865 0.9 ;
			RECT 6.775 0.43 7.005 0.9 ;
			RECT 5.915 0.43 6.145 0.9 ;
			RECT 5.915 0.43 7.865 0.66 ;
			RECT 6.345 3.1 7.435 3.33 ;
			RECT 7.205 0.89 7.435 3.33 ;
			RECT 6.345 2.665 6.575 3.33 ;
			RECT 1.435 3.375 3.905 3.605 ;
			RECT 3.675 2.505 3.905 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 2.725 2.945 2.955 3.235 ;
			RECT 1.865 2.945 2.095 3.235 ;
			RECT 1.865 3.005 2.955 3.175 ;
			RECT 8.155 0.68 8.385 3.45 ;
			RECT 4.965 1.145 5.195 2.795 ;
			RECT 4.535 0.705 4.765 3.235 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 3.245 0.705 3.475 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFRX4

MACRO ADDFX1
	CLASS CORE ;
	FOREIGN ADDFX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.82 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN CO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 6.31 2.52 6.575 3.53 ;
			RECT 6.31 0.61 6.575 1.26 ;
			RECT 6.31 0.61 6.57 3.53 ;

		END 

	END CO
	PIN S
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 7.205 2.52 7.49 3.53 ;
			RECT 7.23 0.61 7.49 3.53 ;
			RECT 7.205 0.61 7.49 1.26 ;

		END 

	END S
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.745 3.81 2.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.41587 LAYER met1  ;
		ANTENNAMAXAREACAR 1.34111 LAYER met1  ;
		ANTENNAGATEAREA 0.63 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 0.955 4.73 2.195 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.41587 LAYER met1  ;
		ANTENNAMAXAREACAR 1.34111 LAYER met1  ;
		ANTENNAGATEAREA 0.63 LAYER met1  ;
	END B
	PIN CI
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.47 4.27 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.88783 LAYER met1  ;
		ANTENNAMAXAREACAR 1.72698 LAYER met1  ;
		ANTENNAGATEAREA 0.4725 LAYER met1  ;
	END CI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.82 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.82 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.825 0.6 6.055 0.89 ;
			RECT 3.675 0.6 3.905 0.89 ;
			RECT 2.815 0.6 3.045 0.89 ;
			RECT 2.815 0.675 6.055 0.815 ;
			RECT 5.395 2.59 5.625 2.88 ;
			RECT 5.44 1.125 5.58 2.88 ;
			RECT 5.395 1.125 5.625 1.415 ;
			RECT 2.295 0.655 2.525 0.945 ;
			RECT 1.435 0.655 1.665 0.945 ;
			RECT 1.435 0.73 2.525 0.87 ;
			RECT 0.975 3.15 1.265 3.32 ;
			RECT 1.05 0.655 1.19 3.32 ;
			RECT 1.005 2.0 1.235 2.29 ;
			RECT 1.005 0.655 1.235 0.945 ;
			RECT 2.785 3.15 6.085 3.32 ;
			RECT 1.405 3.15 2.555 3.32 ;

	END

END ADDFX1

MACRO AOI22X1
	CLASS CORE ;
	FOREIGN AOI22X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.435 2.82 1.97 3.11 ;
			RECT 1.71 0.82 1.97 3.11 ;
			RECT 0.975 0.82 1.97 1.05 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.83 0.59 2.07 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.24 1.05 2.48 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.525573 LAYER met1  ;
		ANTENNAMAXAREACAR 0.446737 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.195 2.43 2.435 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.699824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.596085 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.205 1.51 2.445 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.546737 LAYER met1  ;
		ANTENNAMAXAREACAR 0.464727 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 3.3 2.125 3.53 ;
			RECT 1.005 2.88 1.235 3.53 ;
			RECT 0.145 2.88 0.375 3.53 ;

	END

END AOI22X1

MACRO SDFFRX4
	CLASS CORE ;
	FOREIGN SDFFRX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 14.72 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 12.115 0.68 12.55 3.45 ;
			RECT 11.255 1.77 12.55 2.0 ;
			RECT 11.255 0.68 11.485 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 13.835 0.675 14.065 3.45 ;
			RECT 13.67 0.675 14.065 3.445 ;
			RECT 12.975 1.77 14.065 2.0 ;
			RECT 12.975 0.68 13.205 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.4 2.43 1.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.13 1.05 3.37 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.17 5.19 2.41 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.48112 LAYER met1  ;
		ANTENNAMAXAREACAR 1.39499 LAYER met1  ;
		ANTENNAGATEAREA 0.609 LAYER met1  ;
	END RN
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.16508 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08206 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.78 2.43 3.02 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 14.72 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 14.72 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 9.445 0.88 9.675 3.315 ;
			RECT 8.585 2.665 8.815 3.315 ;
			RECT 8.585 2.665 9.675 2.895 ;
			RECT 8.115 2.195 9.675 2.425 ;
			RECT 6.775 0.705 7.005 3.235 ;
			RECT 6.775 1.855 7.545 2.085 ;
			RECT 3.675 3.375 6.145 3.605 ;
			RECT 5.915 2.475 6.145 3.605 ;
			RECT 3.675 0.705 3.905 3.605 ;
			RECT 1.435 3.375 3.475 3.605 ;
			RECT 3.245 0.705 3.475 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 10.395 0.68 10.625 3.45 ;
			RECT 8.125 0.57 10.135 0.74 ;
			RECT 7.715 1.145 7.945 2.795 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.485 0.705 5.715 3.235 ;
			RECT 4.075 3.005 5.225 3.175 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFRX4

MACRO CLKBUFX8
	CLASS CORE ;
	FOREIGN CLKBUFX8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.06 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 0.68 4.27 3.45 ;
			RECT 1.435 2.44 4.27 2.67 ;
			RECT 1.435 0.68 4.27 0.91 ;
			RECT 3.155 2.44 3.385 3.45 ;
			RECT 3.155 0.68 3.385 1.33 ;
			RECT 2.295 2.44 2.525 3.45 ;
			RECT 2.295 0.68 2.525 1.33 ;
			RECT 1.435 2.44 1.665 3.45 ;
			RECT 1.435 0.68 1.665 1.33 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.415 0.59 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.336861 LAYER met1  ;
		ANTENNAMAXAREACAR 0.337302 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.06 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.06 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 3.235 1.02 3.525 ;
			RECT 0.73 0.61 1.02 3.525 ;
			RECT 0.73 1.51 1.57 1.74 ;
			RECT 0.575 0.61 1.02 0.9 ;

	END

END CLKBUFX8

MACRO AOI21X1
	CLASS CORE ;
	FOREIGN AOI21X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.435 2.635 1.97 2.925 ;
			RECT 1.71 0.61 1.97 2.925 ;
			RECT 1.005 0.61 1.97 0.9 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 0.0007 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.00023 LAYER met1  ;
	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.775 0.59 2.015 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.447972 LAYER met1  ;
		ANTENNAMAXAREACAR 0.380776 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.685 1.05 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.409171 LAYER met1  ;
		ANTENNAMAXAREACAR 0.347795 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.04 1.51 2.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.44515 LAYER met1  ;
		ANTENNAMAXAREACAR 0.378995 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.265 3.5 ;

	END

END AOI21X1

MACRO OAI221X2
	CLASS CORE ;
	FOREIGN OAI221X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.98 BY 4.135 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.435 2.87 5.65 3.1 ;
			RECT 5.39 1.48 5.65 3.1 ;
			RECT 5.055 1.48 5.65 1.71 ;
			RECT 5.055 2.87 5.285 3.52 ;
			RECT 5.055 1.04 5.285 1.71 ;
			RECT 3.675 2.87 3.905 3.16 ;
			RECT 1.435 2.87 1.665 3.16 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.565 0.59 2.805 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.48 1.51 2.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.485 2.89 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.485 3.81 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 1.465 4.73 2.705 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.439153 LAYER met1  ;
		ANTENNAMAXAREACAR 0.42425 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.98 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.98 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.485 0.61 5.715 1.26 ;
			RECT 4.625 0.61 4.855 1.26 ;
			RECT 3.675 0.61 3.905 0.9 ;
			RECT 2.815 0.61 3.045 0.9 ;
			RECT 2.815 0.61 5.715 0.84 ;
			RECT 0.145 1.1 4.335 1.33 ;
			RECT 4.105 1.04 4.335 1.33 ;
			RECT 3.245 1.04 3.475 1.33 ;
			RECT 2.385 0.68 2.615 1.33 ;
			RECT 1.435 0.68 1.665 1.33 ;
			RECT 0.575 0.68 0.805 1.33 ;
			RECT 2.385 3.3 4.335 3.53 ;
			RECT 4.105 3.24 4.335 3.53 ;
			RECT 3.245 3.24 3.475 3.53 ;
			RECT 2.385 3.24 2.615 3.53 ;
			RECT 0.145 3.3 2.095 3.53 ;
			RECT 1.865 3.24 2.095 3.53 ;
			RECT 1.005 3.23 1.235 3.53 ;
			RECT 0.145 3.23 0.375 3.53 ;

	END

END OAI221X2

MACRO SDFFX4
	CLASS CORE ;
	FOREIGN SDFFX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 12.88 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.365 0.675 10.71 3.45 ;
			RECT 9.505 1.77 10.71 2.0 ;
			RECT 9.505 0.68 9.735 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 12.085 0.675 12.55 3.45 ;
			RECT 11.225 1.77 12.55 2.0 ;
			RECT 11.225 0.68 11.455 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.435 2.43 1.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.15 1.05 3.39 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.745 1.05 1.985 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.16508 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08206 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.82 2.43 3.06 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 12.88 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 12.88 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.675 3.375 5.715 3.605 ;
			RECT 5.485 2.475 5.715 3.605 ;
			RECT 3.675 0.705 3.905 3.605 ;
			RECT 1.435 3.375 3.475 3.605 ;
			RECT 3.245 0.705 3.475 3.605 ;
			RECT 1.435 0.705 1.665 3.605 ;
			RECT 8.645 0.68 8.875 3.45 ;
			RECT 7.695 0.88 7.925 3.315 ;
			RECT 6.775 1.145 7.005 2.795 ;
			RECT 6.345 0.705 6.575 3.235 ;
			RECT 5.915 0.705 6.145 3.235 ;
			RECT 4.965 0.705 5.195 3.235 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFX4

MACRO AOI211X2
	CLASS CORE ;
	FOREIGN AOI211X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 0.7 3.905 3.07 ;
			RECT 1.405 1.035 3.905 1.265 ;
			RECT 2.815 0.97 3.045 1.265 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 0.0007 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.00023 LAYER met1  ;
	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.25 0.59 2.49 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.326279 LAYER met1  ;
		ANTENNAMAXAREACAR 0.328307 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.51 1.51 2.75 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.313933 LAYER met1  ;
		ANTENNAMAXAREACAR 0.317813 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.51 2.89 2.75 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.330864 LAYER met1  ;
		ANTENNAMAXAREACAR 0.34575 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.51 3.35 2.75 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.446208 LAYER met1  ;
		ANTENNAMAXAREACAR 0.430247 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.355 3.26 4.365 3.49 ;
			RECT 0.11 2.89 3.075 3.12 ;
			RECT 0.11 0.64 2.12 0.87 ;

	END

END AOI211X2

MACRO BUFX8
	CLASS CORE ;
	FOREIGN BUFX8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.06 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.435 3.22 4.27 3.51 ;
			RECT 4.01 0.635 4.27 3.51 ;
			RECT 3.155 0.635 3.385 3.51 ;
			RECT 2.295 0.635 2.525 3.51 ;
			RECT 1.435 0.635 1.665 3.51 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.355 0.59 2.595 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.383774 LAYER met1  ;
		ANTENNAMAXAREACAR 0.377178 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.06 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.06 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 2.88 0.805 3.53 ;
			RECT 0.575 2.88 1.26 3.11 ;
			RECT 1.03 0.61 1.26 3.11 ;
			RECT 0.575 0.61 1.26 0.9 ;

	END

END BUFX8

MACRO DLY1X1
	CLASS CORE ;
	FOREIGN DLY1X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.065 0.68 3.35 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.2 1.05 2.44 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.21905 LAYER met1  ;
		ANTENNAMAXAREACAR 1.03619 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;
			RECT 1.865 2.505 2.095 2.795 ;
			RECT 1.865 -0.2 2.005 2.795 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;
			RECT 1.215 1.145 1.445 1.435 ;
			RECT 0.82 2.66 1.355 2.8 ;
			RECT 1.215 1.145 1.355 2.8 ;
			RECT 0.82 2.66 0.96 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.145 2.955 2.375 3.245 ;
			RECT 2.235 0.705 2.375 3.245 ;
			RECT 2.145 1.525 2.375 1.815 ;
			RECT 2.145 0.705 2.375 0.995 ;
			RECT 1.435 2.955 1.725 3.245 ;
			RECT 1.585 0.705 1.725 3.245 ;
			RECT 1.495 1.995 1.725 2.285 ;
			RECT 1.435 0.705 1.725 0.995 ;
			RECT 0.09 2.945 0.375 3.235 ;
			RECT 0.09 0.705 0.26 3.235 ;
			RECT 0.09 1.995 0.375 2.285 ;
			RECT 0.09 0.705 0.375 0.995 ;

	END

END DLY1X1

MACRO CLKINVX8
	CLASS CORE ;
	FOREIGN CLKINVX8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.14 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 3.385 3.53 ;
			RECT 3.09 0.61 3.385 3.53 ;
			RECT 0.575 0.61 3.385 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.165 1.97 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.271605 LAYER met1  ;
		ANTENNAMAXAREACAR 0.307319 LAYER met1  ;
		ANTENNAGATEAREA 2.268 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.14 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.14 4.34 ;

		END 

	END VDD

END CLKINVX8

MACRO NAND4X4
	CLASS CORE ;
	FOREIGN NAND4X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.82 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 7.49 3.53 ;
			RECT 7.23 1.04 7.49 3.53 ;
			RECT 7.115 1.04 7.49 1.33 ;
			RECT 6.255 1.04 6.485 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.43 1.05 2.67 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.45 2.89 2.69 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.44 5.19 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 6.77 1.475 7.03 2.715 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.82 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.82 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.865 0.64 2.095 1.29 ;
			RECT 1.005 0.64 1.235 1.29 ;
			RECT 0.145 0.64 0.375 1.29 ;
			RECT 0.145 0.64 3.845 0.87 ;
			RECT 4.075 0.64 7.805 0.87 ;
			RECT 2.265 1.07 5.655 1.3 ;

	END

END NAND4X4

MACRO NAND2X4
	CLASS CORE ;
	FOREIGN NAND2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.14 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 3.415 3.53 ;
			RECT 3.09 1.07 3.415 3.53 ;
			RECT 2.265 1.07 3.415 1.3 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.36 1.05 2.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.44 2.89 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.14 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.14 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 0.615 3.845 0.905 ;

	END

END NAND2X4

MACRO AND4X1
	CLASS CORE ;
	FOREIGN AND4X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.355 3.24 2.89 3.53 ;
			RECT 2.63 0.61 2.89 3.53 ;
			RECT 2.355 0.61 2.89 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.41 1.97 2.65 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.736508 LAYER met1  ;
		ANTENNAMAXAREACAR 0.626032 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.055 1.51 2.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.725079 LAYER met1  ;
		ANTENNAMAXAREACAR 0.617448 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.89 1.05 3.13 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.657778 LAYER met1  ;
		ANTENNAMAXAREACAR 0.559111 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.055 0.59 2.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.653968 LAYER met1  ;
		ANTENNAMAXAREACAR 0.555873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.545 3.27 2.215 3.5 ;
			RECT 1.985 2.87 2.215 3.5 ;
			RECT 2.17 1.04 2.43 3.1 ;
			RECT 1.985 0.685 2.215 1.27 ;
			RECT 0.115 0.685 2.215 0.915 ;

	END

END AND4X1

MACRO AND2X1
	CLASS CORE ;
	FOREIGN AND2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.495 2.86 1.97 3.51 ;
			RECT 1.71 0.625 1.97 3.51 ;
			RECT 1.495 0.625 1.97 0.915 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.695 0.59 2.935 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.653968 LAYER met1  ;
		ANTENNAMAXAREACAR 0.555873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.155 1.51 2.395 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.2381 LAYER met1  ;
		ANTENNAMAXAREACAR 1.05238 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 3.24 1.11 3.53 ;
			RECT 0.88 0.685 1.11 3.53 ;
			RECT 0.145 0.655 0.375 0.945 ;
			RECT 0.145 0.685 1.11 0.915 ;

	END

END AND2X1

MACRO AOI222X2
	CLASS CORE ;
	FOREIGN AOI222X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.9 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.915 1.04 6.145 3.235 ;
			RECT 5.055 2.945 6.145 3.085 ;
			RECT 5.85 1.04 6.145 3.085 ;
			RECT 1.435 1.04 6.145 1.21 ;
			RECT 5.055 2.945 5.285 3.235 ;
			RECT 3.675 0.92 3.905 1.21 ;
			RECT 1.435 0.92 1.665 1.21 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.24 0.59 2.48 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.333333 LAYER met1  ;
		ANTENNAMAXAREACAR 0.334303 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.42 1.51 2.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.46 2.89 2.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.43 3.81 2.67 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328042 LAYER met1  ;
		ANTENNAMAXAREACAR 0.329806 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.445 5.19 2.685 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.328395 LAYER met1  ;
		ANTENNAMAXAREACAR 0.330388 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 6.31 1.305 6.57 2.545 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.396825 LAYER met1  ;
		ANTENNAMAXAREACAR 0.388272 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.9 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.9 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 6.345 0.61 6.575 0.9 ;
			RECT 5.485 0.61 5.715 0.9 ;
			RECT 4.625 0.61 4.855 0.9 ;
			RECT 4.625 0.61 6.575 0.75 ;
			RECT 2.815 3.405 6.575 3.545 ;
			RECT 6.345 3.255 6.575 3.545 ;
			RECT 5.485 3.255 5.715 3.545 ;
			RECT 4.625 3.255 4.855 3.545 ;
			RECT 3.675 3.255 3.905 3.545 ;
			RECT 2.815 3.255 3.045 3.545 ;
			RECT 4.105 0.61 4.335 0.9 ;
			RECT 3.245 0.61 3.475 0.9 ;
			RECT 2.385 0.61 2.615 0.9 ;
			RECT 2.385 0.61 4.335 0.75 ;
			RECT 4.105 2.945 4.335 3.235 ;
			RECT 3.245 2.945 3.475 3.235 ;
			RECT 2.385 2.945 2.615 3.235 ;
			RECT 1.865 2.945 2.095 3.235 ;
			RECT 1.005 2.945 1.235 3.235 ;
			RECT 0.145 2.945 0.375 3.235 ;
			RECT 0.145 2.945 4.335 3.085 ;
			RECT 1.865 0.61 2.095 0.9 ;
			RECT 1.005 0.61 1.235 0.9 ;
			RECT 0.145 0.61 0.375 0.9 ;
			RECT 0.145 0.61 2.095 0.75 ;

	END

END AOI222X2

MACRO OR3X1
	CLASS CORE ;
	FOREIGN OR3X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.925 3.24 2.43 3.53 ;
			RECT 2.17 0.535 2.43 3.53 ;
			RECT 1.925 0.535 2.43 0.825 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.46 1.51 2.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.692063 LAYER met1  ;
		ANTENNAMAXAREACAR 0.588254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.1 1.05 2.34 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.742857 LAYER met1  ;
		ANTENNAMAXAREACAR 0.631429 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.665 0.59 2.905 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.87 1.2 3.5 ;
			RECT 0.97 2.87 2.03 3.1 ;
			RECT 1.8 1.09 2.03 3.1 ;
			RECT 1.36 1.09 2.03 1.32 ;
			RECT 1.36 0.475 1.59 1.32 ;
			RECT 0.115 0.475 1.59 0.705 ;

	END

END OR3X1

MACRO OAI211X2
	CLASS CORE ;
	FOREIGN OAI211X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 3.035 3.905 3.325 ;
			RECT 3.55 1.04 3.905 1.33 ;
			RECT 1.34 2.805 3.81 3.035 ;
			RECT 3.55 1.04 3.81 3.325 ;
			RECT 2.815 2.805 3.045 3.13 ;
			RECT 1.34 2.805 1.665 3.13 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.415 0.59 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.42 1.51 2.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.41 2.89 2.65 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.48 4.27 2.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.393298 LAYER met1  ;
		ANTENNAMAXAREACAR 0.385273 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.105 0.535 4.335 0.9 ;
			RECT 3.245 0.535 3.475 0.9 ;
			RECT 2.385 0.535 2.615 0.9 ;
			RECT 2.385 0.535 4.335 0.765 ;
			RECT 0.115 1.04 3.075 1.27 ;
			RECT 0.115 3.27 2.125 3.5 ;

	END

END OAI211X2

MACRO INVX8
	CLASS CORE ;
	FOREIGN INVX8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.14 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 3.385 3.53 ;
			RECT 3.09 0.675 3.385 3.53 ;
			RECT 0.575 0.675 3.385 0.965 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.315 1.05 2.555 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.313051 LAYER met1  ;
		ANTENNAMAXAREACAR 0.355291 LAYER met1  ;
		ANTENNAGATEAREA 2.268 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.14 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.14 4.34 ;

		END 

	END VDD

END INVX8

MACRO AOI221X2
	CLASS CORE ;
	FOREIGN AOI221X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.98 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.05 2.43 5.715 2.69 ;
			RECT 5.39 0.59 5.715 2.69 ;
			RECT 4.62 0.59 5.715 0.85 ;
			RECT 5.05 2.43 5.31 3.08 ;
			RECT 1.435 1.05 4.88 1.19 ;
			RECT 4.62 0.59 4.88 1.19 ;
			RECT 3.675 0.9 3.905 1.19 ;
			RECT 1.435 0.9 1.665 1.19 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.19 0.59 2.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.389771 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382275 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.4 1.51 2.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.389771 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382275 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.415 3.35 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.234568 LAYER met1  ;
		ANTENNAMAXAREACAR 0.199383 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.42 2.43 2.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.213404 LAYER met1  ;
		ANTENNAMAXAREACAR 0.181393 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 1.425 4.73 2.665 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.439153 LAYER met1  ;
		ANTENNAMAXAREACAR 0.42425 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.98 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.98 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.265 3.24 5.745 3.41 ;
			RECT 2.355 0.59 4.365 0.76 ;
			RECT 0.115 2.88 3.845 3.05 ;
			RECT 0.115 0.59 2.125 0.76 ;

	END

END AOI221X2

MACRO TBUFX1
	CLASS CORE ;
	FOREIGN TBUFX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 3.09 2.52 3.535 3.53 ;
			RECT 3.09 0.61 3.535 1.26 ;
			RECT 3.09 0.61 3.35 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.665 1.97 2.905 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.911111 LAYER met1  ;
		ANTENNAMAXAREACAR 0.86619 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END A
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.85 1.05 3.09 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.50476 LAYER met1  ;
		ANTENNAMAXAREACAR 1.37079 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END OE
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.385 3.24 2.615 3.53 ;
			RECT 2.43 0.785 2.57 3.53 ;
			RECT 2.385 1.82 2.615 2.11 ;
			RECT 2.375 0.785 2.605 1.075 ;
			RECT 1.435 3.24 1.665 3.53 ;
			RECT 1.43 0.685 1.57 3.385 ;
			RECT 1.34 1.48 1.57 1.77 ;
			RECT 1.005 0.61 1.235 0.9 ;
			RECT 1.005 0.685 1.62 0.825 ;
			RECT 0.145 3.24 0.375 3.53 ;
			RECT 0.175 0.61 0.345 3.53 ;
			RECT 0.145 1.82 0.375 2.11 ;
			RECT 0.145 0.61 0.375 0.9 ;

	END

END TBUFX1

MACRO SDFFSRX4
	CLASS CORE ;
	FOREIGN SDFFSRX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 17.02 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 14.59 0.68 14.935 3.45 ;
			RECT 13.735 1.77 14.935 2.0 ;
			RECT 13.735 0.68 13.965 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 16.315 0.68 16.69 3.455 ;
			RECT 15.455 1.77 16.69 2.0 ;
			RECT 15.455 0.68 15.685 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 2.02 2.43 3.26 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.13651 LAYER met1  ;
		ANTENNAMAXAREACAR 0.966032 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.36 1.05 3.6 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.679365 LAYER met1  ;
		ANTENNAMAXAREACAR 0.57746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.145 3.81 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END RN
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.945 1.05 2.185 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.08571 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0146 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.635 2.43 1.875 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.780952 LAYER met1  ;
		ANTENNAMAXAREACAR 0.66381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.56 3.39 11.545 3.59 ;
			RECT 11.345 2.245 11.545 3.59 ;
			RECT 11.16 2.245 11.545 2.535 ;
			RECT 5.56 1.145 5.79 3.59 ;
			RECT 5.39 1.145 5.79 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.10476 LAYER met1  ;
		ANTENNAMAXAREACAR 0.939048 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 17.02 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 17.02 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 8.155 2.945 8.475 3.235 ;
			RECT 8.245 0.705 8.475 3.235 ;
			RECT 5.02 2.945 5.285 3.235 ;
			RECT 5.02 0.705 5.25 3.235 ;
			RECT 5.02 0.705 5.285 0.995 ;
			RECT 3.18 2.945 3.475 3.235 ;
			RECT 3.18 0.705 3.41 3.235 ;
			RECT 3.18 0.705 3.475 0.995 ;
			RECT 12.875 0.68 13.105 3.45 ;
			RECT 11.925 0.88 12.155 3.315 ;
			RECT 10.115 0.995 11.265 1.165 ;
			RECT 9.595 3.005 11.175 3.175 ;
			RECT 9.595 0.57 10.835 0.74 ;
			RECT 9.195 0.705 9.425 3.235 ;
			RECT 8.765 0.705 8.995 3.235 ;
			RECT 5.975 0.57 7.125 0.74 ;
			RECT 6.435 1.145 6.665 3.235 ;
			RECT 4.625 0.705 4.855 3.235 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFSRX4

MACRO ADDHX1
	CLASS CORE ;
	FOREIGN ADDHX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.06 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN CO
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 2.44 4.885 3.09 ;
			RECT 4.47 0.68 4.885 1.33 ;
			RECT 4.47 0.68 4.73 3.09 ;

		END 

	END CO
	PIN S
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.145 2.44 0.59 3.09 ;
			RECT 0.33 0.68 0.59 3.09 ;
			RECT 0.145 0.68 0.59 1.33 ;

		END 

	END S
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.425 2.43 2.665 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.46667 LAYER met1  ;
		ANTENNAMAXAREACAR 1.33841 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.84 3.81 3.08 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.998942 LAYER met1  ;
		ANTENNAMAXAREACAR 0.984974 LAYER met1  ;
		ANTENNAGATEAREA 0.4725 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.06 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.06 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.735 3.22 4.18 3.51 ;
			RECT 3.95 1.46 4.18 3.51 ;
			RECT 3.305 1.46 4.18 1.69 ;
			RECT 3.305 0.705 3.535 1.69 ;
			RECT 0.73 3.63 2.155 3.8 ;
			RECT 1.895 2.89 2.155 3.8 ;
			RECT 0.73 2.0 0.9 3.8 ;
			RECT 1.605 2.89 2.155 3.06 ;
			RECT 1.605 1.115 1.775 3.06 ;
			RECT 0.73 2.0 1.08 2.29 ;
			RECT 1.605 1.115 2.155 1.285 ;
			RECT 1.925 0.705 2.155 1.285 ;
			RECT 1.22 3.2 1.725 3.49 ;
			RECT 1.22 0.615 1.45 3.49 ;
			RECT 1.22 0.615 1.725 0.905 ;
			RECT 2.785 0.705 3.015 3.235 ;

	END

END ADDHX1

MACRO MX4X4
	CLASS CORE ;
	FOREIGN MX4X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 8.74 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 7.635 0.68 7.95 3.45 ;
			RECT 6.775 1.77 7.95 2.0 ;
			RECT 6.775 0.68 7.005 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.85 1.05 3.09 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 2.39 2.43 3.63 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.19 0.905 2.45 2.145 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.02222 LAYER met1  ;
		ANTENNAMAXAREACAR 0.868889 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 2.19 3.81 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.20635 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN S0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.725 1.145 2.955 2.815 ;
			RECT 1.25 1.145 1.51 3.01 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 1.4875 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.4849 LAYER met1  ;
		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 6.44415 LAYER met1  ;
		ANTENNAMAXAREACAR 3.82784 LAYER met1  ;
		ANTENNAGATEAREA 0.4725 LAYER met1  ;
	END S0
	PIN S1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 0.925 4.27 2.165 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.324263 LAYER met1  ;
		ANTENNAMAXAREACAR 0.341156 LAYER met1  ;
		ANTENNAGATEAREA 0.441 LAYER met1  ;
	END S1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 8.74 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 8.74 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.155 3.57 6.055 3.8 ;
			RECT 5.825 0.68 6.055 3.8 ;
			RECT 3.155 0.705 3.385 3.8 ;
			RECT 1.435 3.24 1.88 3.53 ;
			RECT 1.65 0.61 1.88 3.53 ;
			RECT 1.435 0.61 1.88 0.9 ;
			RECT 5.395 0.68 5.625 3.235 ;
			RECT 4.965 0.68 5.195 3.235 ;
			RECT 4.445 0.705 4.675 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END MX4X4

MACRO MX2X4
	CLASS CORE ;
	FOREIGN MX2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.845 3.235 4.27 3.525 ;
			RECT 4.01 0.61 4.27 3.525 ;
			RECT 2.845 0.61 4.27 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.175 1.05 2.415 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.469546 LAYER met1  ;
		ANTENNAMAXAREACAR 0.399114 LAYER met1  ;
		ANTENNAGATEAREA 0.22575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.255 3.35 2.495 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.2979 LAYER met1  ;
		ANTENNAMAXAREACAR 1.10321 LAYER met1  ;
		ANTENNAGATEAREA 0.22575 LAYER met1  ;
	END B
	PIN S0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.405 1.51 2.645 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.887149 LAYER met1  ;
		ANTENNAMAXAREACAR 0.862161 LAYER met1  ;
		ANTENNAGATEAREA 0.38325 LAYER met1  ;
	END S0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.495 3.025 2.235 3.315 ;
			RECT 2.005 1.025 2.235 3.315 ;
			RECT 2.005 2.03 2.47 2.26 ;
			RECT 1.495 1.025 2.235 1.255 ;
			RECT 1.495 0.705 1.725 1.255 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END MX2X4

MACRO OAI21X1
	CLASS CORE ;
	FOREIGN OAI21X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.005 3.24 1.97 3.53 ;
			RECT 1.71 0.61 1.97 3.53 ;
			RECT 1.435 0.61 1.97 0.9 ;
			RECT 1.005 2.795 1.235 3.53 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.165 0.59 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.325 1.05 2.565 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.245 1.51 2.485 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.536155 LAYER met1  ;
		ANTENNAMAXAREACAR 0.455732 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 0.64 1.265 0.87 ;

	END

END OAI21X1

MACRO DFFSRX1
	CLASS CORE ;
	FOREIGN DFFSRX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 11.5 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.245 2.42 10.71 3.57 ;
			RECT 10.45 0.57 10.71 3.57 ;
			RECT 10.245 0.57 10.71 1.35 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 10.91 2.42 11.275 3.57 ;
			RECT 10.91 0.57 11.275 1.35 ;
			RECT 10.91 0.57 11.17 3.57 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.1873 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00921 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.805 1.05 2.045 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.742857 LAYER met1  ;
		ANTENNAMAXAREACAR 0.631429 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 6.77 1.155 7.03 2.395 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.02222 LAYER met1  ;
		ANTENNAMAXAREACAR 0.868889 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END RN
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.075 4.27 2.315 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.95238 LAYER met1  ;
		ANTENNAMAXAREACAR 1.75127 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 11.5 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 11.5 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.945 0.845 8.545 1.015 ;
			RECT 8.315 0.705 8.545 1.015 ;
			RECT 5.945 0.705 6.175 1.015 ;
			RECT 5.555 3.425 8.545 3.595 ;
			RECT 8.315 3.26 8.545 3.595 ;
			RECT 5.555 3.26 5.785 3.595 ;
			RECT 5.125 2.535 5.355 3.235 ;
			RECT 5.125 2.535 8.38 2.765 ;
			RECT 5.515 0.705 5.745 2.765 ;
			RECT 7.885 2.945 8.115 3.235 ;
			RECT 6.415 2.945 6.645 3.235 ;
			RECT 6.415 3.005 8.115 3.175 ;
			RECT 3.405 3.005 4.925 3.235 ;
			RECT 4.695 0.715 4.925 3.235 ;
			RECT 3.405 2.945 3.635 3.235 ;
			RECT 4.695 0.715 5.315 0.945 ;
			RECT 5.085 0.655 5.315 0.945 ;
			RECT 1.435 3.405 3.265 3.575 ;
			RECT 3.095 2.165 3.265 3.575 ;
			RECT 1.435 0.705 1.665 3.575 ;
			RECT 3.095 2.165 3.325 2.455 ;
			RECT 9.695 0.705 9.925 3.235 ;
			RECT 8.835 0.705 9.065 3.235 ;
			RECT 6.345 0.535 8.145 0.705 ;
			RECT 3.215 0.715 4.365 0.885 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFSRX1

MACRO CLKINVX1
	CLASS CORE ;
	FOREIGN CLKINVX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.545 2.905 1.05 3.495 ;
			RECT 0.79 0.64 1.05 3.495 ;
			RECT 0.545 0.64 1.05 0.87 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.19 0.59 2.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD

END CLKINVX1

MACRO NOR4X2
	CLASS CORE ;
	FOREIGN NOR4X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 2.83 3.905 3.12 ;
			RECT 0.545 0.61 3.905 0.9 ;
			RECT 3.55 0.61 3.81 3.12 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.205 0.59 2.445 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.415 1.51 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.205 2.89 2.445 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.299824 LAYER met1  ;
		ANTENNAMAXAREACAR 0.30582 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.44 4.27 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.393298 LAYER met1  ;
		ANTENNAMAXAREACAR 0.385273 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.355 3.27 4.365 3.5 ;
			RECT 1.405 2.9 3.075 3.13 ;
			RECT 0.115 3.27 2.125 3.5 ;

	END

END NOR4X2

MACRO NOR2X2
	CLASS CORE ;
	FOREIGN NOR2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 2.445 1.665 3.095 ;
			RECT 1.25 0.68 1.665 1.33 ;
			RECT 1.25 0.68 1.51 3.095 ;
			RECT 0.575 0.68 1.665 0.94 ;
			RECT 0.575 0.68 0.805 1.33 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.49 0.59 2.73 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.319224 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32231 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.49 2.43 2.73 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.502646 LAYER met1  ;
		ANTENNAMAXAREACAR 0.478219 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.11 3.27 2.125 3.5 ;

	END

END NOR2X2

MACRO NAND3X1
	CLASS CORE ;
	FOREIGN NAND3X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.16 1.97 3.45 ;
			RECT 1.71 0.61 1.97 3.45 ;
			RECT 1.435 0.61 1.97 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.165 0.59 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.497354 LAYER met1  ;
		ANTENNAMAXAREACAR 0.422751 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.685 1.05 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.47 1.51 2.71 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.546737 LAYER met1  ;
		ANTENNAMAXAREACAR 0.464727 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD

END NAND3X1

MACRO XOR2X2
	CLASS CORE ;
	FOREIGN XOR2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.77 3.2 3.35 3.495 ;
			RECT 3.09 0.605 3.35 3.495 ;
			RECT 2.77 0.605 3.35 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.375 2.43 2.615 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.952381 LAYER met1  ;
		ANTENNAMAXAREACAR 0.809524 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 2.055 0.59 3.295 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.00952 LAYER met1  ;
		ANTENNAMAXAREACAR 1.97794 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 3.32 2.63 3.49 ;
			RECT 2.46 2.875 2.63 3.49 ;
			RECT 2.46 2.875 2.95 3.045 ;
			RECT 2.78 1.065 2.95 3.045 ;
			RECT 2.72 1.485 2.95 1.775 ;
			RECT 2.395 1.065 2.95 1.235 ;
			RECT 2.395 0.535 2.565 1.235 ;
			RECT 1.405 0.535 2.565 0.705 ;
			RECT 1.025 2.98 2.125 3.15 ;
			RECT 1.025 0.845 1.285 3.15 ;
			RECT 1.025 0.845 2.125 1.015 ;
			RECT 0.01 3.44 0.375 3.73 ;
			RECT 0.01 0.655 0.18 3.73 ;
			RECT 0.01 1.61 0.375 1.9 ;
			RECT 0.01 0.655 0.375 0.945 ;

	END

END XOR2X2

MACRO INVX1
	CLASS CORE ;
	FOREIGN INVX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 2.84 1.05 3.49 ;
			RECT 0.79 0.605 1.05 3.49 ;
			RECT 0.575 0.605 1.05 1.255 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.43 0.59 2.67 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD

END INVX1

MACRO XNOR2X1
	CLASS CORE ;
	FOREIGN XNOR2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.77 2.44 3.35 2.7 ;
			RECT 3.09 1.055 3.35 2.7 ;
			RECT 2.77 1.055 3.35 1.315 ;
			RECT 2.77 2.44 3.03 3.09 ;
			RECT 2.77 0.61 3.03 1.315 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.435 1.05 2.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.730159 LAYER met1  ;
		ANTENNAMAXAREACAR 0.620635 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.87 0.59 2.11 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.99365 LAYER met1  ;
		ANTENNAMAXAREACAR 2.05619 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.365 1.665 3.655 ;
			RECT 1.435 3.365 2.63 3.595 ;
			RECT 2.46 0.64 2.63 3.595 ;
			RECT 2.4 1.49 2.63 1.78 ;
			RECT 1.405 0.64 2.63 0.87 ;
			RECT 1.005 2.975 1.235 3.655 ;
			RECT 1.005 2.975 1.67 3.145 ;
			RECT 1.5 1.105 1.67 3.145 ;
			RECT 1.5 2.03 2.27 2.26 ;
			RECT 1.005 1.105 1.67 1.275 ;
			RECT 1.005 0.64 1.235 1.275 ;
			RECT 0.015 3.24 0.375 3.53 ;
			RECT 0.015 0.39 0.185 3.53 ;
			RECT 0.015 2.385 0.295 2.675 ;
			RECT 0.015 0.39 0.375 0.68 ;

	END

END XNOR2X1

MACRO TBUFX8
	CLASS CORE ;
	FOREIGN TBUFX8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 9.2 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 8.125 0.68 8.41 3.45 ;
			RECT 5.545 1.58 8.41 1.81 ;
			RECT 7.265 0.68 7.495 3.45 ;
			RECT 6.405 0.68 6.635 3.45 ;
			RECT 5.545 0.68 5.775 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.04 1.97 2.28 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.5 LAYER met1  ;
		ANTENNAMAXAREACAR 0.501455 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.57 3.625 3.8 ;
			RECT 3.395 1.98 3.625 3.8 ;
			RECT 0.575 2.97 0.805 3.8 ;
			RECT 0.33 1.98 0.59 3.22 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.7245 LAYER met1  ;
	END OE
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 9.2 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 9.2 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.825 3.345 6.205 3.575 ;
			RECT 5.975 2.0 6.205 3.575 ;
			RECT 4.685 1.12 4.915 3.575 ;
			RECT 3.825 2.42 4.055 3.575 ;
			RECT 4.165 1.12 4.915 1.35 ;
			RECT 4.165 0.945 4.395 1.35 ;
			RECT 2.445 2.8 2.675 3.09 ;
			RECT 2.445 2.8 3.12 3.0 ;
			RECT 2.92 1.525 3.12 3.0 ;
			RECT 5.115 0.555 5.345 1.77 ;
			RECT 2.34 1.525 3.12 1.725 ;
			RECT 2.34 0.555 2.54 1.725 ;
			RECT 1.065 0.555 1.295 1.33 ;
			RECT 1.925 0.555 2.155 0.9 ;
			RECT 1.065 0.555 5.345 0.785 ;
			RECT 2.785 1.125 3.965 1.355 ;
			RECT 3.735 0.945 3.965 1.355 ;
			RECT 2.785 0.945 3.015 1.355 ;
			RECT 1.065 3.23 3.105 3.43 ;
			RECT 2.875 3.14 3.105 3.43 ;
			RECT 2.015 3.14 2.245 3.43 ;
			RECT 1.065 3.14 1.295 3.43 ;
			RECT 0.015 3.39 0.375 3.68 ;
			RECT 0.015 0.705 0.185 3.68 ;
			RECT 1.065 2.425 2.34 2.655 ;
			RECT 2.11 2.03 2.34 2.655 ;
			RECT 1.065 1.51 1.295 2.655 ;
			RECT 2.11 2.03 2.4 2.26 ;
			RECT 0.015 1.51 1.295 1.74 ;
			RECT 0.015 0.705 0.375 0.995 ;

	END

END TBUFX8

MACRO OAI22X1
	CLASS CORE ;
	FOREIGN OAI22X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.975 3.27 2.43 3.5 ;
			RECT 2.17 1.025 2.43 3.5 ;
			RECT 1.405 1.025 2.43 1.255 ;
			RECT 0.975 3.205 1.265 3.5 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.325 1.165 0.585 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.380952 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32381 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.52 1.05 2.76 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.380952 LAYER met1  ;
		ANTENNAMAXAREACAR 0.32381 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.685 1.97 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.409171 LAYER met1  ;
		ANTENNAMAXAREACAR 0.347795 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.42 1.51 2.66 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.398589 LAYER met1  ;
		ANTENNAMAXAREACAR 0.338801 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.835 0.655 2.125 0.885 ;
			RECT 0.975 0.655 1.265 0.885 ;
			RECT 0.115 0.655 0.405 0.885 ;
			RECT 0.115 0.7 2.125 0.84 ;

	END

END OAI22X1

MACRO OR4X1
	CLASS CORE ;
	FOREIGN OR4X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.355 3.24 2.89 3.53 ;
			RECT 2.63 0.535 2.89 3.53 ;
			RECT 2.355 0.535 2.89 0.825 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 0.845 1.51 2.085 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.755556 LAYER met1  ;
		ANTENNAMAXAREACAR 0.642222 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.485 1.97 2.725 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.41905 LAYER met1  ;
		ANTENNAMAXAREACAR 2.32603 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.865 0.59 2.105 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.634921 LAYER met1  ;
		ANTENNAMAXAREACAR 0.539683 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.29 1.05 2.53 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.34286 LAYER met1  ;
		ANTENNAMAXAREACAR 2.26127 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.87 1.2 3.5 ;
			RECT 0.97 2.87 2.37 3.1 ;
			RECT 2.14 1.07 2.37 3.1 ;
			RECT 1.82 1.07 2.37 1.3 ;
			RECT 1.82 0.475 2.05 1.3 ;
			RECT 0.545 0.475 2.05 0.705 ;

	END

END OR4X1

MACRO OR2X1
	CLASS CORE ;
	FOREIGN OR2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.495 3.21 1.97 3.5 ;
			RECT 1.71 0.505 1.97 3.5 ;
			RECT 1.495 0.505 1.97 0.795 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.455 1.05 2.695 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.920635 LAYER met1  ;
		ANTENNAMAXAREACAR 0.78254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.145 0.59 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.27 1.2 3.5 ;
			RECT 0.97 2.84 1.2 3.5 ;
			RECT 1.19 0.965 1.42 3.07 ;
			RECT 0.765 0.965 1.42 1.195 ;
			RECT 0.765 0.475 0.995 1.195 ;
			RECT 0.545 0.475 0.995 0.705 ;

	END

END OR2X1

MACRO BUFX2
	CLASS CORE ;
	FOREIGN BUFX2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.84 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.065 3.23 1.51 3.52 ;
			RECT 1.25 0.61 1.51 3.52 ;
			RECT 1.065 0.61 1.51 1.26 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.685 1.05 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.11746 LAYER met1  ;
		ANTENNAMAXAREACAR 0.949841 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.84 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.84 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 3.24 0.375 3.53 ;
			RECT 0.145 0.655 0.285 3.53 ;
			RECT 0.145 1.48 0.375 1.77 ;
			RECT 0.145 0.655 0.375 0.945 ;

	END

END BUFX2

MACRO XNOR2X4
	CLASS CORE ;
	FOREIGN XNOR2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.52 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.47 2.44 4.885 3.45 ;
			RECT 4.47 0.68 4.885 1.33 ;
			RECT 4.47 0.68 4.73 3.45 ;
			RECT 3.795 1.77 4.73 2.0 ;
			RECT 3.795 0.68 4.025 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 2.085 0.59 3.325 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.005 1.05 2.245 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.478458 LAYER met1  ;
		ANTENNAMAXAREACAR 0.472222 LAYER met1  ;
		ANTENNAGATEAREA 0.441 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.52 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.52 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.985 0.68 2.215 3.09 ;
			RECT 1.985 1.51 3.595 1.74 ;
			RECT 1.525 3.27 3.195 3.5 ;
			RECT 2.905 2.55 3.195 3.5 ;
			RECT 1.525 2.55 1.815 3.5 ;
			RECT 1.615 2.0 1.845 2.29 ;
			RECT 1.615 0.68 1.785 2.29 ;
			RECT 1.555 0.68 1.785 1.33 ;
			RECT 1.005 2.61 1.33 3.235 ;
			RECT 1.19 0.39 1.33 3.235 ;
			RECT 1.19 1.66 1.42 1.95 ;
			RECT 1.005 0.39 1.33 0.865 ;
			RECT 0.01 3.47 0.375 3.76 ;
			RECT 0.01 0.39 0.18 3.76 ;
			RECT 0.01 1.66 0.29 1.95 ;
			RECT 0.01 0.39 0.375 0.68 ;

	END

END XNOR2X4

MACRO INVX4
	CLASS CORE ;
	FOREIGN INVX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 1.695 3.53 ;
			RECT 1.25 0.61 1.695 3.53 ;
			RECT 0.575 0.61 1.695 0.9 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.455 1.05 2.695 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.268078 LAYER met1  ;
		ANTENNAMAXAREACAR 0.304321 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD

END INVX4

MACRO CLKBUFX2
	CLASS CORE ;
	FOREIGN CLKBUFX2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.84 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.065 3.24 1.51 3.53 ;
			RECT 1.25 0.61 1.51 3.53 ;
			RECT 1.065 0.61 1.51 1.26 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.805 1.05 3.045 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.11746 LAYER met1  ;
		ANTENNAMAXAREACAR 0.949841 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 3.24 0.375 3.53 ;
			RECT 0.145 0.655 0.285 3.53 ;
			RECT 0.145 1.48 0.375 1.77 ;
			RECT 0.145 0.655 0.375 0.945 ;

	END

END CLKBUFX2

MACRO CLKAND2X2
	CLASS CORE ;
	FOREIGN CLKAND2X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.49 3.24 1.97 3.53 ;
			RECT 1.71 0.68 1.97 3.53 ;
			RECT 1.495 0.68 1.97 1.33 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.685 1.51 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.845198 LAYER met1  ;
		ANTENNAMAXAREACAR 0.718418 LAYER met1  ;
		ANTENNAGATEAREA 0.22125 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.855 0.59 3.095 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.632768 LAYER met1  ;
		ANTENNAMAXAREACAR 0.537853 LAYER met1  ;
		ANTENNAGATEAREA 0.22125 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 3.24 0.96 3.53 ;
			RECT 0.73 1.55 0.96 3.53 ;

	END

END CLKAND2X2

MACRO DFFSRX4
	CLASS CORE ;
	FOREIGN DFFSRX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 14.72 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 11.83 2.44 12.165 3.45 ;
			RECT 11.83 0.68 12.165 1.33 ;
			RECT 11.83 0.68 12.09 3.45 ;
			RECT 11.075 1.77 12.09 2.0 ;
			RECT 11.075 0.68 11.305 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 13.655 0.68 13.93 3.45 ;
			RECT 12.795 1.77 13.93 2.0 ;
			RECT 12.795 0.68 13.025 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.805 1.05 2.045 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787937 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 6.77 1.62 7.03 2.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.02222 LAYER met1  ;
		ANTENNAMAXAREACAR 0.868889 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END RN
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 4.01 1.06 4.27 2.3 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.94603 LAYER met1  ;
		ANTENNAMAXAREACAR 1.74587 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 14.72 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 14.72 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 5.125 1.25 5.355 3.235 ;
			RECT 8.835 1.25 9.065 2.115 ;
			RECT 5.125 1.25 9.065 1.48 ;
			RECT 5.515 0.705 5.745 1.48 ;
			RECT 5.945 0.88 8.545 1.05 ;
			RECT 8.315 0.705 8.545 1.05 ;
			RECT 5.945 0.705 6.175 1.05 ;
			RECT 5.555 3.405 8.545 3.575 ;
			RECT 8.315 3.24 8.545 3.575 ;
			RECT 5.555 3.24 5.785 3.575 ;
			RECT 7.885 2.945 8.115 3.235 ;
			RECT 6.415 2.945 6.645 3.235 ;
			RECT 6.415 3.005 8.115 3.175 ;
			RECT 3.405 3.005 4.925 3.235 ;
			RECT 4.695 0.715 4.925 3.235 ;
			RECT 3.405 2.945 3.635 3.235 ;
			RECT 4.695 0.715 5.315 0.945 ;
			RECT 5.085 0.655 5.315 0.945 ;
			RECT 1.435 3.405 3.265 3.575 ;
			RECT 3.095 2.165 3.265 3.575 ;
			RECT 1.435 0.705 1.665 3.575 ;
			RECT 3.095 2.165 3.325 2.455 ;
			RECT 10.215 0.68 10.445 3.45 ;
			RECT 9.265 0.88 9.495 3.315 ;
			RECT 6.345 0.57 8.145 0.74 ;
			RECT 3.215 0.57 4.365 0.74 ;
			RECT 2.725 0.705 2.955 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DFFSRX4

MACRO CLKINVX4
	CLASS CORE ;
	FOREIGN CLKINVX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.3 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 1.97 3.53 ;
			RECT 1.71 0.64 1.97 3.53 ;
			RECT 0.575 0.64 1.97 0.93 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.455 0.59 2.695 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.097884 LAYER met1  ;
		ANTENNAMAXAREACAR 0.083201 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.3 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.3 4.34 ;

		END 

	END VDD

END CLKINVX4

MACRO NAND3X4
	CLASS CORE ;
	FOREIGN NAND3X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.44 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.24 6.11 3.53 ;
			RECT 5.85 0.65 6.11 3.53 ;
			RECT 4.075 1.07 6.11 1.3 ;
			RECT 5.825 0.65 6.11 1.3 ;
			RECT 4.075 1.07 4.305 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.48 1.05 2.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.44 2.89 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.93 1.44 5.19 2.68 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.239859 LAYER met1  ;
		ANTENNAMAXAREACAR 0.25485 LAYER met1  ;
		ANTENNAGATEAREA 1.134 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.44 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.44 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.145 1.07 3.845 1.3 ;
			RECT 1.865 0.65 2.095 1.3 ;
			RECT 1.005 0.65 1.235 1.3 ;
			RECT 0.145 0.65 0.375 1.3 ;
			RECT 2.265 0.64 5.655 0.87 ;

	END

END NAND3X4

MACRO AND3X1
	CLASS CORE ;
	FOREIGN AND3X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.385 3.045 2.89 3.335 ;
			RECT 2.63 0.69 2.89 3.335 ;
			RECT 2.385 0.69 2.89 0.98 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 0.815 0.59 2.055 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.890159 LAYER met1  ;
		ANTENNAMAXAREACAR 0.756635 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.705 1.05 2.945 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.933333 LAYER met1  ;
		ANTENNAMAXAREACAR 0.793333 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.03 1.51 2.27 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.661587 LAYER met1  ;
		ANTENNAMAXAREACAR 0.562349 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.005 3.175 1.235 3.465 ;
			RECT 0.145 3.175 0.375 3.465 ;
			RECT 0.145 3.175 2.19 3.405 ;
			RECT 1.96 0.64 2.19 3.405 ;
			RECT 1.405 0.64 2.19 0.87 ;

	END

END AND3X1

MACRO AOI211X1
	CLASS CORE ;
	FOREIGN AOI211X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.87 2.79 2.43 3.08 ;
			RECT 2.17 0.64 2.43 3.08 ;
			RECT 0.115 0.64 2.43 0.87 ;
			RECT 0.115 0.64 0.405 1.23 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 0.0007 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.00023 LAYER met1  ;
	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.05 1.05 2.29 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.57 0.59 2.81 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.363316 LAYER met1  ;
		ANTENNAMAXAREACAR 0.308818 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.57 1.51 2.81 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.38448 LAYER met1  ;
		ANTENNAMAXAREACAR 0.326808 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.29 1.97 2.53 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.405644 LAYER met1  ;
		ANTENNAMAXAREACAR 0.344797 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.005 3.18 1.235 3.47 ;
			RECT 0.145 3.18 0.375 3.47 ;
			RECT 0.145 3.21 1.235 3.44 ;

	END

END AOI211X1

MACRO OAI221X1
	CLASS CORE ;
	FOREIGN OAI221X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.815 0.61 3.045 1.555 ;
			RECT 0.975 3.27 2.89 3.5 ;
			RECT 2.265 3.025 2.89 3.5 ;
			RECT 2.63 1.325 2.89 3.5 ;
			RECT 0.975 3.025 1.265 3.5 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.395 0.59 2.635 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.412698 LAYER met1  ;
		ANTENNAMAXAREACAR 0.350794 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.4 1.05 2.64 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.430335 LAYER met1  ;
		ANTENNAMAXAREACAR 0.365785 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.415 1.97 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.43739 LAYER met1  ;
		ANTENNAMAXAREACAR 0.371781 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.225 1.405 1.485 2.645 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.37037 LAYER met1  ;
		ANTENNAMAXAREACAR 0.314815 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.415 2.43 2.655 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.433862 LAYER met1  ;
		ANTENNAMAXAREACAR 0.368783 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.385 0.655 2.615 0.945 ;
			RECT 1.405 0.685 1.695 0.915 ;
			RECT 1.405 0.73 2.615 0.87 ;
			RECT 1.835 1.025 2.125 1.255 ;
			RECT 0.975 1.025 1.265 1.255 ;
			RECT 0.115 1.025 0.405 1.255 ;
			RECT 0.115 1.07 2.125 1.21 ;

	END

END OAI221X1

MACRO SDFFSRX1
	CLASS CORE ;
	FOREIGN SDFFSRX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 14.72 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 13.23 0.68 13.575 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 14.13 0.675 14.425 3.45 ;

		END 

	END QN
	PIN CK
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 2.17 2.02 2.43 3.26 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.13651 LAYER met1  ;
		ANTENNAMAXAREACAR 0.966032 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.785 2.46 1.05 3.7 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.907937 LAYER met1  ;
		ANTENNAMAXAREACAR 0.771746 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.145 3.81 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END RN
	PIN SE
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.945 1.05 2.185 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.08571 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0146 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SE
	PIN SI
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.635 2.43 1.875 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.780952 LAYER met1  ;
		ANTENNAMAXAREACAR 0.66381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SI
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.425 3.39 11.545 3.59 ;
			RECT 11.345 2.245 11.545 3.59 ;
			RECT 11.16 2.245 11.545 2.535 ;
			RECT 5.425 1.15 5.685 3.75 ;
			RECT 5.39 1.145 5.65 2.385 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.10476 LAYER met1  ;
		ANTENNAMAXAREACAR 0.939048 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 14.72 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 14.72 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 8.155 2.945 8.475 3.235 ;
			RECT 8.245 0.705 8.475 3.235 ;
			RECT 5.02 2.945 5.285 3.235 ;
			RECT 5.02 0.705 5.25 3.235 ;
			RECT 5.02 0.705 5.285 0.995 ;
			RECT 3.095 2.945 3.475 3.235 ;
			RECT 3.095 0.705 3.325 3.235 ;
			RECT 3.095 0.705 3.475 0.995 ;
			RECT 2.57 2.945 2.955 3.235 ;
			RECT 2.57 0.705 2.8 3.235 ;
			RECT 2.57 1.485 2.915 1.775 ;
			RECT 2.57 0.705 2.955 0.995 ;
			RECT 12.815 0.705 13.045 3.235 ;
			RECT 11.865 0.705 12.095 3.235 ;
			RECT 10.115 0.995 11.265 1.165 ;
			RECT 9.595 3.005 11.175 3.175 ;
			RECT 9.595 0.57 10.835 0.74 ;
			RECT 9.195 0.705 9.425 3.235 ;
			RECT 8.765 0.705 8.995 3.235 ;
			RECT 5.975 0.57 7.125 0.74 ;
			RECT 6.435 1.145 6.665 3.235 ;
			RECT 4.625 0.705 4.855 3.235 ;
			RECT 4.105 0.705 4.335 3.235 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END SDFFSRX1

MACRO TBUFX4
	CLASS CORE ;
	FOREIGN TBUFX4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 5.06 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 4.165 0.68 4.73 3.45 ;
			RECT 3.305 1.06 4.73 1.29 ;
			RECT 3.305 0.68 3.535 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.995 1.05 3.235 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.746032 LAYER met1  ;
		ANTENNAMAXAREACAR 0.787037 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN OE
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.925 0.34 2.155 1.77 ;
			RECT 0.575 0.34 2.155 0.57 ;
			RECT 0.575 0.34 0.805 1.79 ;
			RECT 0.33 1.425 0.59 2.665 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.926984 LAYER met1  ;
		ANTENNAMAXAREACAR 0.818519 LAYER met1  ;
		ANTENNAGATEAREA 0.441 LAYER met1  ;
	END OE
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 5.06 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 5.06 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.525 3.345 4.025 3.575 ;
			RECT 3.795 1.46 4.025 3.575 ;
			RECT 1.955 1.91 2.185 3.575 ;
			RECT 1.525 3.24 1.695 3.575 ;
			RECT 1.555 1.91 2.185 2.14 ;
			RECT 1.555 0.71 1.785 2.14 ;
			RECT 1.035 0.71 1.785 0.94 ;
			RECT 2.445 1.525 2.675 3.09 ;
			RECT 2.445 2.03 3.135 2.26 ;
			RECT 2.355 0.68 2.585 1.755 ;
			RECT 0.015 3.63 1.385 3.8 ;
			RECT 1.215 1.49 1.385 3.8 ;
			RECT 0.015 3.24 0.375 3.8 ;
			RECT 0.015 0.705 0.185 3.8 ;
			RECT 1.075 1.48 1.305 1.77 ;
			RECT 0.015 0.705 0.375 0.995 ;

	END

END TBUFX4

MACRO MX4X1
	CLASS CORE ;
	FOREIGN MX4X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.36 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 6.77 0.68 7.03 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.85 1.05 3.09 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.920635 LAYER met1  ;
		ANTENNAMAXAREACAR 0.78254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 2.435 2.43 3.675 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04127 LAYER met1  ;
		ANTENNAMAXAREACAR 0.885079 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.005 2.43 2.245 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.04762 LAYER met1  ;
		ANTENNAMAXAREACAR 0.890476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.815 3.81 3.055 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.20635 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN S0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.725 1.145 2.955 2.815 ;
			RECT 1.25 1.15 1.51 3.065 ;

		END 

		ANTENNAPARTIALMETALSIDEAREA 1.5225 LAYER met1  ;
		ANTENNAPARTIALMETALAREA 0.4979 LAYER met1  ;
		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 6.51822 LAYER met1  ;
		ANTENNAMAXAREACAR 3.85536 LAYER met1  ;
		ANTENNAGATEAREA 0.4725 LAYER met1  ;
	END S0
	PIN S1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 4.01 0.895 4.27 2.135 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.457143 LAYER met1  ;
		ANTENNAMAXAREACAR 0.480317 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END S1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.36 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.36 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 3.155 3.375 6.055 3.605 ;
			RECT 5.825 0.68 6.055 3.605 ;
			RECT 3.155 0.705 3.385 3.605 ;
			RECT 1.435 3.24 1.88 3.53 ;
			RECT 1.65 0.705 1.88 3.53 ;
			RECT 1.435 0.705 1.88 0.995 ;
			RECT 5.395 0.68 5.625 3.235 ;
			RECT 4.965 0.68 5.195 3.235 ;
			RECT 4.445 0.705 4.675 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END MX4X1

MACRO MX2X1
	CLASS CORE ;
	FOREIGN MX2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.755 2.91 3.35 3.5 ;
			RECT 3.09 0.64 3.35 3.5 ;
			RECT 2.755 0.64 3.35 1.23 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.48 1.05 1.72 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.653968 LAYER met1  ;
		ANTENNAMAXAREACAR 0.555873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 0.875 2.43 2.115 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.793651 LAYER met1  ;
		ANTENNAMAXAREACAR 0.674603 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END B
	PIN S0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.28 1.05 3.52 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.06032 LAYER met1  ;
		ANTENNAMAXAREACAR 2.11286 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END S0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 0.655 1.665 3.38 ;
			RECT 1.435 2.29 2.84 2.52 ;
			RECT 2.61 2.0 2.84 2.52 ;
			RECT 0.145 0.655 0.375 3.38 ;

	END

END MX2X1

MACRO DLY4X4
	CLASS CORE ;
	FOREIGN DLY4X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 11.5 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 10.395 0.68 10.71 3.45 ;
			RECT 9.535 1.77 10.71 2.0 ;
			RECT 9.535 0.68 9.765 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.20635 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 11.505 0.2 ;
			RECT 5.395 -0.2 5.625 2.815 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 11.5 4.34 ;
			RECT 3.155 1.125 3.385 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 8.675 0.68 8.905 3.235 ;
			RECT 8.155 0.705 8.385 3.235 ;
			RECT 6.435 0.705 6.665 3.235 ;
			RECT 5.915 0.705 6.145 3.235 ;
			RECT 4.195 0.705 4.425 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 1.955 0.705 2.185 3.235 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DLY4X4

MACRO DLY2X4
	CLASS CORE ;
	FOREIGN DLY2X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.9 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.85 0.68 6.145 3.45 ;
			RECT 5.055 1.77 6.145 2.0 ;
			RECT 5.055 0.68 5.285 3.45 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.19 1.05 3.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.20635 LAYER met1  ;
		ANTENNAMAXAREACAR 1.0254 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.905 0.2 ;
			RECT 2.6 -0.2 2.83 2.815 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.905 4.34 ;
			RECT 3.155 1.125 3.385 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.195 0.68 4.425 3.235 ;
			RECT 3.675 0.705 3.905 3.235 ;
			RECT 1.955 0.705 2.185 3.235 ;
			RECT 1.435 0.705 1.665 3.235 ;
			RECT 0.145 0.705 0.375 3.235 ;

	END

END DLY2X4

MACRO AOI21X2
	CLASS CORE ;
	FOREIGN AOI21X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.215 0.625 3.505 1.23 ;
			RECT 0.575 0.625 3.505 0.915 ;
			RECT 0.575 2.755 1.05 3.045 ;
			RECT 0.79 0.625 1.05 3.045 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.565 1.51 2.805 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.296296 LAYER met1  ;
		ANTENNAMAXAREACAR 0.302822 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.56 2.89 2.8 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.296296 LAYER met1  ;
		ANTENNAMAXAREACAR 0.302822 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.27 0.59 2.51 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.301587 LAYER met1  ;
		ANTENNAMAXAREACAR 0.307319 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.115 3.24 3.505 3.47 ;
			RECT 1.405 1.07 3.07 1.3 ;

	END

END AOI21X2

MACRO CLKXOR2X1
	CLASS CORE ;
	FOREIGN CLKXOR2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.22 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 0.62 2.985 3.495 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.595 1.05 2.835 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.653968 LAYER met1  ;
		ANTENNAMAXAREACAR 0.555873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.925 0.59 3.165 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 2.00952 LAYER met1  ;
		ANTENNAMAXAREACAR 1.97794 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.22 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.22 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.405 3.32 2.49 3.49 ;
			RECT 2.23 0.535 2.49 3.49 ;
			RECT 1.405 0.535 2.49 0.705 ;
			RECT 0.975 2.98 1.995 3.15 ;
			RECT 1.735 0.845 1.995 3.15 ;
			RECT 0.975 0.845 1.995 1.015 ;
			RECT 0.02 3.38 0.405 3.55 ;
			RECT 0.02 0.655 0.19 3.55 ;
			RECT 0.02 1.495 0.3 1.785 ;
			RECT 0.02 0.655 0.375 0.945 ;

	END

END CLKXOR2X1

MACRO DLY1X4
	CLASS CORE ;
	FOREIGN DLY1X4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.815 3.36 3.905 3.53 ;
			RECT 3.55 0.61 3.905 3.53 ;
			RECT 2.815 0.61 3.905 0.84 ;
			RECT 2.815 0.61 3.045 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.62 1.05 1.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.27619 LAYER met1  ;
		ANTENNAMAXAREACAR 1.08476 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END A
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;
			RECT 1.095 2.505 1.36 2.795 ;
			RECT 1.19 -0.2 1.36 2.795 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;
			RECT 0.725 2.0 0.955 2.29 ;
			RECT 0.755 2.0 0.925 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.955 3.24 2.185 3.53 ;
			RECT 1.985 0.61 2.155 3.53 ;
			RECT 1.955 2.0 2.185 2.29 ;
			RECT 1.955 0.61 2.185 0.9 ;
			RECT 1.435 3.24 1.665 3.53 ;
			RECT 1.5 0.61 1.67 3.385 ;
			RECT 1.5 1.485 1.73 1.775 ;
			RECT 1.5 0.61 1.73 0.9 ;
			RECT 0.145 3.24 0.375 3.53 ;
			RECT 0.175 0.61 0.345 3.53 ;
			RECT 0.14 1.485 0.37 1.775 ;
			RECT 0.145 0.61 0.375 0.9 ;

	END

END DLY1X4

MACRO AOI22X2
	CLASS CORE ;
	FOREIGN AOI22X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 4.6 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.815 2.95 4.27 3.09 ;
			RECT 4.01 1.05 4.27 3.09 ;
			RECT 1.435 1.05 4.27 1.19 ;
			RECT 3.675 2.95 3.905 3.24 ;
			RECT 2.815 2.95 3.045 3.24 ;
			RECT 2.815 0.9 3.045 1.19 ;
			RECT 1.435 0.9 1.665 1.19 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.52 0.59 2.76 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.389771 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382275 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.39 1.51 2.63 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.389771 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382275 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.55 1.355 3.81 2.595 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.390123 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382857 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.52 2.89 2.76 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.389771 LAYER met1  ;
		ANTENNAMAXAREACAR 0.382275 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 4.6 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 4.6 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 2.355 0.59 4.365 0.76 ;
			RECT 0.115 3.38 4.365 3.55 ;
			RECT 0.115 0.59 2.125 0.76 ;

	END

END AOI22X2

MACRO NOR3X2
	CLASS CORE ;
	FOREIGN NOR3X2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 2.8 3.045 3.09 ;
			RECT 0.575 0.61 3.045 0.9 ;
			RECT 2.63 0.61 2.89 3.09 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.33 0.59 2.57 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.405644 LAYER met1  ;
		ANTENNAMAXAREACAR 0.395767 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.455 1.97 2.695 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.405644 LAYER met1  ;
		ANTENNAMAXAREACAR 0.395767 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.295 3.35 2.535 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.322751 LAYER met1  ;
		ANTENNAMAXAREACAR 0.325309 LAYER met1  ;
		ANTENNAGATEAREA 0.567 LAYER met1  ;
	END C
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.495 3.27 3.505 3.5 ;
			RECT 0.545 2.9 2.215 3.13 ;

	END

END NOR3X2

MACRO NAND4X1
	CLASS CORE ;
	FOREIGN NAND4X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 2.76 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.23 2.43 3.52 ;
			RECT 2.17 0.61 2.43 3.52 ;
			RECT 1.865 0.61 2.43 0.9 ;
			RECT 1.435 3.23 1.665 3.53 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.685 0.59 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.511464 LAYER met1  ;
		ANTENNAMAXAREACAR 0.434744 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.165 1.05 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.514991 LAYER met1  ;
		ANTENNAMAXAREACAR 0.437743 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN C
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.685 1.51 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.536155 LAYER met1  ;
		ANTENNAMAXAREACAR 0.455732 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C
	PIN D
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.165 1.97 2.405 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.557319 LAYER met1  ;
		ANTENNAMAXAREACAR 0.473721 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END D
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 2.76 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 2.76 4.34 ;

		END 

	END VDD

END NAND4X1

MACRO NAND2X1
	CLASS CORE ;
	FOREIGN NAND2X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.84 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 3.21 1.51 3.47 ;
			RECT 1.25 0.655 1.51 3.47 ;
			RECT 0.975 0.655 1.51 0.915 ;
			RECT 0.575 2.82 0.805 3.47 ;

		END 

	END Y
	PIN A
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.29 0.59 2.53 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.504409 LAYER met1  ;
		ANTENNAMAXAREACAR 0.428748 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A
	PIN B
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.19 1.05 2.43 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.514991 LAYER met1  ;
		ANTENNAMAXAREACAR 0.437743 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.84 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.84 4.34 ;

		END 

	END VDD

END NAND2X1

MACRO OAI222X1
	CLASS CORE ;
	FOREIGN OAI222X1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.63 1.04 3.045 1.33 ;
			RECT 1.005 3.3 2.89 3.53 ;
			RECT 2.63 1.04 2.89 3.53 ;
			RECT 2.385 3.24 2.89 3.53 ;
			RECT 1.005 3.24 1.235 3.53 ;

		END 

	END Y
	PIN A0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.33 1.38 0.59 2.62 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.493827 LAYER met1  ;
		ANTENNAMAXAREACAR 0.419753 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A0
	PIN A1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 1.685 1.05 2.925 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.493827 LAYER met1  ;
		ANTENNAMAXAREACAR 0.419753 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END A1
	PIN B0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.25 1.39 1.51 2.63 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.645503 LAYER met1  ;
		ANTENNAMAXAREACAR 0.548677 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B0
	PIN B1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 1.71 1.58 1.97 2.82 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.673721 LAYER met1  ;
		ANTENNAMAXAREACAR 0.572663 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END B1
	PIN C0
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 3.09 1.62 3.35 2.86 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.47619 LAYER met1  ;
		ANTENNAMAXAREACAR 0.404762 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C0
	PIN C1
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 2.17 1.385 2.43 2.625 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.652557 LAYER met1  ;
		ANTENNAMAXAREACAR 0.554674 LAYER met1  ;
		ANTENNAGATEAREA 0.2835 LAYER met1  ;
	END C1
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.495 0.64 3.505 0.87 ;
			RECT 0.545 1.01 2.215 1.24 ;

	END

END OAI222X1

MACRO FILL1
	CLASS CORE ;
	FOREIGN FILL1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.46 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 0.46 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 0.46 4.34 ;

		END 

	END VDD

END FILL1

MACRO FILL2
	CLASS CORE ;
	FOREIGN FILL2 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 0.92 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 0.92 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 0.92 4.34 ;

		END 

	END VDD

END FILL2

MACRO FILL4
	CLASS CORE ;
	FOREIGN FILL4 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.84 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.84 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.84 4.34 ;

		END 

	END VDD

END FILL4

MACRO FILL8
	CLASS CORE ;
	FOREIGN FILL8 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 3.68 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 3.68 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 3.68 4.34 ;

		END 

	END VDD

END FILL8

MACRO FILL16
	CLASS CORE ;
	FOREIGN FILL16 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 7.36 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 7.36 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 7.36 4.34 ;

		END 

	END VDD

END FILL16

MACRO FILL32
	CLASS CORE ;
	FOREIGN FILL32 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 14.72 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 14.72 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 14.72 4.34 ;

		END 

	END VDD

END FILL32

MACRO FILL64
	CLASS CORE ;
	FOREIGN FILL64 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 29.44 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 29.44 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 29.44 4.34 ;

		END 

	END VDD

END FILL64

MACRO TIEHI
	CLASS CORE ;
	FOREIGN TIEHI 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.575 2.84 1.05 3.49 ;
			RECT 0.79 2.25 1.05 3.49 ;

		END 

	END Y
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 0.575 0.605 0.805 1.255 ;

	END

END TIEHI

MACRO TIELO
	CLASS CORE ;
	FOREIGN TIELO 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 1.38 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Y
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.605 1.05 1.845 ;
			RECT 0.575 0.605 1.05 1.255 ;

		END 

	END Y
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 1.38 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		SHAPE ABUTMENT ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 1.38 4.34 ;

		END 

	END VDD

END TIELO

MACRO TLATX1
	CLASS CORE ;
	FOREIGN TLATX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.9 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.39 0.68 5.65 3.45 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 6.275 2.44 6.57 3.45 ;
			RECT 6.31 0.68 6.57 3.45 ;
			RECT 6.275 0.68 6.57 1.33 ;

		END 

	END QN
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.34 1.05 3.255 ;
			RECT 0.735 2.505 1.05 2.795 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.05397 LAYER met1  ;
		ANTENNAMAXAREACAR 0.895873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN G
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.83 1.05 1.75 ;
			RECT 0.72 1.145 1.05 1.435 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END G
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.9 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.9 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 1.435 3.485 3.46 3.715 ;
			RECT 3.23 0.415 3.46 3.715 ;
			RECT 1.435 2.945 1.665 3.715 ;
			RECT 1.435 0.415 1.665 0.995 ;
			RECT 1.435 0.415 3.46 0.645 ;
			RECT 2.645 2.505 2.875 2.795 ;
			RECT 2.7 1.145 2.84 2.795 ;
			RECT 2.645 1.145 2.875 1.435 ;
			RECT 4.665 0.68 4.895 3.45 ;
			RECT 3.715 0.705 3.945 3.235 ;
			RECT 0.075 0.705 0.305 3.235 ;

	END

END TLATX1

MACRO TLATSRX1
	CLASS CORE ;
	FOREIGN TLATSRX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 8.74 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN Q
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 7.09 2.44 7.49 3.45 ;
			RECT 7.23 0.68 7.49 3.45 ;
			RECT 7.09 0.68 7.49 1.33 ;

		END 

	END Q
	PIN QN
		DIRECTION OUTPUT ;
		PORT 
			LAYER met1 ;
			RECT 7.95 2.44 8.41 3.45 ;
			RECT 8.15 0.68 8.41 3.45 ;
			RECT 7.95 0.68 8.41 1.33 ;

		END 

	END QN
	PIN D
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 1.25 2.34 1.51 3.255 ;
			RECT 1.165 2.505 1.51 2.795 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.05397 LAYER met1  ;
		ANTENNAMAXAREACAR 0.895873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END D
	PIN G
		DIRECTION INPUT ;
		USE CLOCK ;
		PORT 
			LAYER met1 ;
			RECT 0.33 2.34 0.59 3.255 ;
			RECT 0.12 2.34 0.59 2.57 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 0.634921 LAYER met1  ;
		ANTENNAMAXAREACAR 0.539683 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END G
	PIN RN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 1.24 0.815 3.86 0.955 ;
			RECT 3.57 0.725 3.86 0.955 ;
			RECT 3.55 0.815 3.81 1.77 ;
			RECT 1.15 1.145 1.38 1.435 ;
			RECT 1.24 0.815 1.38 1.435 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.315 LAYER met1  ;
	END RN
	PIN SN
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 5.39 1.43 5.65 2.205 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.50476 LAYER met1  ;
		ANTENNAMAXAREACAR 1.27905 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END SN
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS!" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 8.74 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD!" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 8.74 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.96 2.945 5.19 3.235 ;
			RECT 4.96 3.02 6.2 3.16 ;
			RECT 6.06 1.485 6.2 3.16 ;
			RECT 5.97 1.485 6.2 1.775 ;
			RECT 1.91 3.66 4.82 3.8 ;
			RECT 4.68 2.57 4.82 3.8 ;
			RECT 1.91 2.945 2.05 3.8 ;
			RECT 1.865 2.945 2.095 3.235 ;
			RECT 4.68 2.57 5.465 2.71 ;
			RECT 5.05 2.42 5.465 2.71 ;
			RECT 5.05 0.34 5.19 2.71 ;
			RECT 1.865 0.34 2.095 0.63 ;
			RECT 1.865 0.34 5.19 0.48 ;
			RECT 4.18 2.185 4.41 2.475 ;
			RECT 4.215 1.145 4.355 2.475 ;
			RECT 4.18 1.145 4.41 1.435 ;
			RECT 6.34 0.68 6.57 3.45 ;

	END

END TLATSRX1

MACRO ICGX1
	CLASS CORE ;
	FOREIGN ICGX1 0.0 0.0  ;
	ORIGIN 0.0 0.0 ;
	SIZE 6.44 BY 4.14 ;
	SYMMETRY X Y ;
	SITE CoreSite ;
	PIN ECK
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT 
			LAYER met1 ;
			RECT 5.85 2.86 6.12 3.51 ;
			RECT 5.85 0.625 6.11 3.51 ;
			RECT 5.82 0.61 6.05 0.9 ;

		END 

	END ECK
	PIN CK
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 0.83 1.05 1.75 ;
			RECT 0.72 1.145 1.05 1.435 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.18095 LAYER met1  ;
		ANTENNAMAXAREACAR 1.00381 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END CK
	PIN E
		DIRECTION INPUT ;
		PORT 
			LAYER met1 ;
			RECT 0.79 2.34 1.05 3.255 ;

		END 

		ANTENNAMODEL OXIDE1 ;
		ANTENNAMAXSIDEAREACAR 1.05397 LAYER met1  ;
		ANTENNAMAXAREACAR 0.895873 LAYER met1  ;
		ANTENNAGATEAREA 0.1575 LAYER met1  ;
	END E
	PIN VSS
		DIRECTION INPUT ;
		USE GROUND ;
		NETEXPR "VSS VSS" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 -0.2 6.44 0.2 ;

		END 

	END VSS
	PIN VDD
		DIRECTION INPUT ;
		USE POWER ;
		NETEXPR "VDD VDD" ;
		PORT 
			LAYER met1 ;
			RECT 0.0 3.94 6.44 4.34 ;

		END 

	END VDD
	OBS
			LAYER met1 ;
			RECT 4.985 0.685 5.215 3.46 ;
			RECT 4.485 0.655 4.715 0.945 ;
			RECT 4.485 0.685 5.215 0.915 ;
			RECT 1.435 3.485 3.46 3.715 ;
			RECT 3.23 0.415 3.46 3.715 ;
			RECT 1.435 2.945 1.665 3.715 ;
			RECT 1.435 0.415 1.665 0.995 ;
			RECT 1.435 0.415 3.46 0.645 ;
			RECT 2.645 2.505 2.875 2.795 ;
			RECT 2.7 1.145 2.84 2.795 ;
			RECT 2.645 1.145 2.875 1.435 ;
			RECT 3.715 0.705 3.945 3.235 ;
			RECT 0.145 0.695 0.375 3.235 ;

	END

END ICGX1

END LIBRARY
